
module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n66, n67, n69, n70, n73,
         n74, n75, n76, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n128,
         n129, n131, n132, n134, n135, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n216, n219, n221, n222, n223, n224, n225, n226, n227, n229, n230,
         n231, n232, n233, n234, n235, n236, n244, n274, n275, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n346, n347, n348, n349, n350, n351, n352, n353;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U103 ( .A(n145), .B(n151), .CI(n100), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n153), .B(n166), .CI(n159), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n170), .B(n163), .CO(n123), .S(n124) );
  BUF_X1 U237 ( .A(n234), .Z(n304) );
  BUF_X1 U238 ( .A(n236), .Z(n295) );
  BUF_X2 U239 ( .A(n216), .Z(n286) );
  INV_X1 U240 ( .A(n320), .ZN(n66) );
  CLKBUF_X1 U241 ( .A(n50), .Z(n274) );
  OR2_X1 U242 ( .A1(n118), .A2(n121), .ZN(n275) );
  AND3_X1 U243 ( .A1(n279), .A2(n280), .A3(n281), .ZN(product[15]) );
  OR2_X1 U244 ( .A1(n172), .A2(n140), .ZN(n277) );
  XOR2_X1 U245 ( .A(n141), .B(n83), .Z(n278) );
  XOR2_X1 U246 ( .A(n14), .B(n278), .Z(product[14]) );
  NAND2_X1 U247 ( .A1(n14), .A2(n141), .ZN(n279) );
  NAND2_X1 U248 ( .A1(n14), .A2(n83), .ZN(n280) );
  NAND2_X1 U249 ( .A1(n141), .A2(n83), .ZN(n281) );
  OR2_X2 U250 ( .A1(n307), .A2(n306), .ZN(n283) );
  XNOR2_X1 U251 ( .A(n282), .B(n120), .ZN(n118) );
  XNOR2_X1 U252 ( .A(n161), .B(n168), .ZN(n282) );
  BUF_X2 U253 ( .A(n235), .Z(n346) );
  OR2_X1 U254 ( .A1(n307), .A2(n306), .ZN(n221) );
  BUF_X1 U255 ( .A(n225), .Z(n349) );
  INV_X1 U256 ( .A(n229), .ZN(n284) );
  OR2_X2 U257 ( .A1(n305), .A2(n135), .ZN(n288) );
  AOI21_X1 U258 ( .B1(n343), .B2(n67), .A(n320), .ZN(n62) );
  BUF_X2 U259 ( .A(n348), .Z(n285) );
  BUF_X2 U260 ( .A(n235), .Z(n348) );
  XNOR2_X1 U261 ( .A(n310), .B(n131), .ZN(n94) );
  NAND2_X1 U262 ( .A1(n226), .A2(n339), .ZN(n287) );
  OR2_X1 U263 ( .A1(n305), .A2(n135), .ZN(n224) );
  XNOR2_X1 U264 ( .A(n295), .B(a[2]), .ZN(n289) );
  NOR2_X1 U265 ( .A1(n101), .A2(n96), .ZN(n35) );
  BUF_X1 U266 ( .A(n97), .Z(n290) );
  CLKBUF_X1 U267 ( .A(n234), .Z(n291) );
  XNOR2_X2 U268 ( .A(n346), .B(a[4]), .ZN(n292) );
  CLKBUF_X1 U269 ( .A(n236), .Z(n293) );
  CLKBUF_X1 U270 ( .A(n236), .Z(n294) );
  BUF_X2 U271 ( .A(n289), .Z(n296) );
  BUF_X1 U272 ( .A(n227), .Z(n350) );
  XOR2_X1 U273 ( .A(n119), .B(n154), .Z(n297) );
  XOR2_X1 U274 ( .A(n116), .B(n297), .Z(n114) );
  NAND2_X1 U275 ( .A1(n116), .A2(n119), .ZN(n298) );
  NAND2_X1 U276 ( .A1(n116), .A2(n154), .ZN(n299) );
  NAND2_X1 U277 ( .A1(n119), .A2(n154), .ZN(n300) );
  NAND3_X1 U278 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n113) );
  CLKBUF_X1 U279 ( .A(n44), .Z(n301) );
  NOR2_X1 U280 ( .A1(n113), .A2(n108), .ZN(n44) );
  XNOR2_X1 U281 ( .A(n302), .B(n94), .ZN(n92) );
  XNOR2_X1 U282 ( .A(n97), .B(n144), .ZN(n302) );
  CLKBUF_X1 U283 ( .A(n47), .Z(n303) );
  XNOR2_X1 U284 ( .A(n295), .B(n135), .ZN(n305) );
  INV_X1 U285 ( .A(n135), .ZN(n244) );
  XNOR2_X1 U286 ( .A(a[6]), .B(n233), .ZN(n306) );
  XOR2_X1 U287 ( .A(n234), .B(a[6]), .Z(n307) );
  CLKBUF_X1 U288 ( .A(n36), .Z(n308) );
  CLKBUF_X1 U289 ( .A(n45), .Z(n309) );
  XOR2_X1 U290 ( .A(n150), .B(n99), .Z(n310) );
  NAND2_X1 U291 ( .A1(n150), .A2(n99), .ZN(n311) );
  NAND2_X1 U292 ( .A1(n150), .A2(n157), .ZN(n312) );
  NAND2_X1 U293 ( .A1(n99), .A2(n157), .ZN(n313) );
  NAND3_X1 U294 ( .A1(n311), .A2(n312), .A3(n313), .ZN(n93) );
  NAND2_X1 U295 ( .A1(n290), .A2(n144), .ZN(n314) );
  NAND2_X1 U296 ( .A1(n290), .A2(n94), .ZN(n315) );
  NAND2_X1 U297 ( .A1(n144), .A2(n94), .ZN(n316) );
  NAND3_X1 U298 ( .A1(n314), .A2(n315), .A3(n316), .ZN(n91) );
  XOR2_X1 U299 ( .A(n348), .B(a[2]), .Z(n317) );
  XNOR2_X1 U300 ( .A(n104), .B(n318), .ZN(n102) );
  XNOR2_X1 U301 ( .A(n109), .B(n106), .ZN(n318) );
  OR2_X1 U302 ( .A1(n114), .A2(n117), .ZN(n319) );
  AND2_X1 U303 ( .A1(n171), .A2(n164), .ZN(n320) );
  NOR2_X1 U304 ( .A1(n35), .A2(n322), .ZN(n321) );
  CLKBUF_X1 U305 ( .A(n324), .Z(n322) );
  AOI21_X1 U306 ( .B1(n55), .B2(n275), .A(n52), .ZN(n50) );
  XNOR2_X1 U307 ( .A(n323), .B(n98), .ZN(n96) );
  XNOR2_X1 U308 ( .A(n103), .B(n105), .ZN(n323) );
  NOR2_X1 U309 ( .A1(n92), .A2(n95), .ZN(n324) );
  NAND2_X1 U310 ( .A1(n219), .A2(n289), .ZN(n325) );
  NAND2_X1 U311 ( .A1(n227), .A2(n317), .ZN(n326) );
  NOR2_X1 U312 ( .A1(n92), .A2(n95), .ZN(n30) );
  NAND2_X1 U313 ( .A1(n289), .A2(n219), .ZN(n223) );
  NAND2_X1 U314 ( .A1(n98), .A2(n103), .ZN(n327) );
  NAND2_X1 U315 ( .A1(n98), .A2(n105), .ZN(n328) );
  NAND2_X1 U316 ( .A1(n103), .A2(n105), .ZN(n329) );
  NAND3_X1 U317 ( .A1(n327), .A2(n328), .A3(n329), .ZN(n95) );
  OAI22_X1 U318 ( .A1(n326), .A2(n192), .B1(n191), .B2(n350), .ZN(n330) );
  NAND2_X1 U319 ( .A1(n120), .A2(n161), .ZN(n331) );
  NAND2_X1 U320 ( .A1(n120), .A2(n168), .ZN(n332) );
  NAND2_X1 U321 ( .A1(n161), .A2(n168), .ZN(n333) );
  NAND3_X1 U322 ( .A1(n331), .A2(n332), .A3(n333), .ZN(n117) );
  NAND2_X1 U323 ( .A1(n226), .A2(n339), .ZN(n334) );
  NAND2_X1 U324 ( .A1(n339), .A2(n226), .ZN(n222) );
  NAND2_X1 U325 ( .A1(n104), .A2(n109), .ZN(n335) );
  NAND2_X1 U326 ( .A1(n104), .A2(n106), .ZN(n336) );
  NAND2_X1 U327 ( .A1(n109), .A2(n106), .ZN(n337) );
  NAND3_X1 U328 ( .A1(n335), .A2(n336), .A3(n337), .ZN(n101) );
  AOI21_X1 U329 ( .B1(n39), .B2(n303), .A(n40), .ZN(n338) );
  OR2_X1 U330 ( .A1(n88), .A2(n91), .ZN(n342) );
  XOR2_X1 U331 ( .A(n234), .B(a[4]), .Z(n339) );
  NOR2_X1 U332 ( .A1(n102), .A2(n107), .ZN(n340) );
  XNOR2_X1 U333 ( .A(n37), .B(n4), .ZN(product[9]) );
  INV_X1 U334 ( .A(n35), .ZN(n74) );
  XOR2_X1 U335 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U336 ( .A1(n342), .A2(n26), .ZN(n2) );
  INV_X1 U337 ( .A(n26), .ZN(n24) );
  OAI21_X1 U338 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  NOR2_X1 U339 ( .A1(n102), .A2(n107), .ZN(n41) );
  INV_X1 U340 ( .A(n19), .ZN(n17) );
  NAND2_X1 U341 ( .A1(n275), .A2(n54), .ZN(n8) );
  NAND2_X1 U342 ( .A1(n344), .A2(n19), .ZN(n1) );
  XOR2_X1 U343 ( .A(n10), .B(n62), .Z(product[3]) );
  INV_X1 U344 ( .A(n60), .ZN(n80) );
  XOR2_X1 U345 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U346 ( .A1(n73), .A2(n31), .ZN(n3) );
  AOI21_X1 U347 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U348 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U349 ( .A1(n76), .A2(n309), .ZN(n6) );
  INV_X1 U350 ( .A(n301), .ZN(n76) );
  XNOR2_X1 U351 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U352 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U353 ( .B1(n46), .B2(n301), .A(n309), .ZN(n43) );
  INV_X1 U354 ( .A(n59), .ZN(n58) );
  XNOR2_X1 U355 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U356 ( .A1(n343), .A2(n66), .ZN(n11) );
  XOR2_X1 U357 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U358 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U359 ( .A(n56), .ZN(n79) );
  NAND2_X1 U360 ( .A1(n319), .A2(n49), .ZN(n7) );
  INV_X1 U361 ( .A(n54), .ZN(n52) );
  OR2_X1 U362 ( .A1(n158), .A2(n146), .ZN(n105) );
  NOR2_X1 U363 ( .A1(n124), .A2(n139), .ZN(n60) );
  XNOR2_X1 U364 ( .A(n70), .B(n341), .ZN(product[13]) );
  XNOR2_X1 U365 ( .A(n85), .B(n84), .ZN(n341) );
  XNOR2_X1 U366 ( .A(n158), .B(n146), .ZN(n106) );
  NOR2_X1 U367 ( .A1(n122), .A2(n123), .ZN(n56) );
  NAND2_X1 U368 ( .A1(n108), .A2(n113), .ZN(n45) );
  NOR2_X1 U369 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U370 ( .A(n83), .ZN(n84) );
  OR2_X1 U371 ( .A1(n171), .A2(n164), .ZN(n343) );
  NAND2_X1 U372 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U373 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U374 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U375 ( .A1(n122), .A2(n123), .ZN(n57) );
  NAND2_X1 U376 ( .A1(n92), .A2(n95), .ZN(n31) );
  OR2_X1 U377 ( .A1(n87), .A2(n86), .ZN(n344) );
  AND2_X1 U378 ( .A1(n286), .A2(n132), .ZN(n164) );
  OR2_X1 U379 ( .A1(n286), .A2(n231), .ZN(n199) );
  INV_X1 U380 ( .A(n128), .ZN(n149) );
  INV_X1 U381 ( .A(n89), .ZN(n90) );
  AND2_X1 U382 ( .A1(n286), .A2(n129), .ZN(n156) );
  OR2_X1 U383 ( .A1(n286), .A2(n230), .ZN(n190) );
  AND2_X1 U384 ( .A1(n277), .A2(n69), .ZN(product[1]) );
  INV_X1 U385 ( .A(n134), .ZN(n165) );
  AND2_X1 U386 ( .A1(n286), .A2(n307), .ZN(n148) );
  INV_X1 U387 ( .A(n125), .ZN(n141) );
  INV_X1 U388 ( .A(n330), .ZN(n100) );
  OR2_X1 U389 ( .A1(n216), .A2(n229), .ZN(n181) );
  OR2_X1 U390 ( .A1(n286), .A2(n232), .ZN(n208) );
  AND2_X1 U391 ( .A1(n286), .A2(n135), .ZN(product[0]) );
  CLKBUF_X1 U392 ( .A(n235), .Z(n347) );
  XNOR2_X1 U393 ( .A(n284), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U394 ( .A(n284), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U395 ( .A(n284), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U396 ( .A(n216), .B(n233), .ZN(n180) );
  INV_X1 U397 ( .A(n233), .ZN(n229) );
  XNOR2_X1 U398 ( .A(n234), .B(a[6]), .ZN(n225) );
  XNOR2_X1 U399 ( .A(n346), .B(a[4]), .ZN(n226) );
  XNOR2_X1 U400 ( .A(n295), .B(a[2]), .ZN(n227) );
  INV_X1 U401 ( .A(n308), .ZN(n34) );
  NAND2_X1 U402 ( .A1(n74), .A2(n308), .ZN(n4) );
  XNOR2_X1 U403 ( .A(n284), .B(b[6]), .ZN(n174) );
  OAI21_X1 U404 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  NAND2_X1 U405 ( .A1(n80), .A2(n61), .ZN(n10) );
  NAND2_X1 U406 ( .A1(n124), .A2(n139), .ZN(n61) );
  INV_X1 U407 ( .A(n131), .ZN(n157) );
  XNOR2_X1 U408 ( .A(n233), .B(b[7]), .ZN(n173) );
  NAND2_X1 U409 ( .A1(n70), .A2(n85), .ZN(n351) );
  NAND2_X1 U410 ( .A1(n70), .A2(n84), .ZN(n352) );
  NAND2_X1 U411 ( .A1(n85), .A2(n84), .ZN(n353) );
  NAND3_X1 U412 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n14) );
  NAND2_X1 U413 ( .A1(n118), .A2(n121), .ZN(n54) );
  INV_X1 U414 ( .A(n347), .ZN(n231) );
  XNOR2_X1 U415 ( .A(n285), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U416 ( .A(n347), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U417 ( .A(n347), .B(b[5]), .ZN(n193) );
  OAI22_X1 U418 ( .A1(n288), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  NAND2_X1 U419 ( .A1(n172), .A2(n140), .ZN(n69) );
  OAI22_X1 U420 ( .A1(n288), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U421 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U422 ( .A1(n288), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U423 ( .A1(n288), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI22_X1 U424 ( .A1(n288), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  OAI22_X1 U425 ( .A1(n224), .A2(n200), .B1(n244), .B2(n200), .ZN(n134) );
  OAI22_X1 U426 ( .A1(n288), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  NAND2_X1 U427 ( .A1(n96), .A2(n101), .ZN(n36) );
  INV_X1 U428 ( .A(n69), .ZN(n67) );
  OAI22_X1 U429 ( .A1(n288), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  XOR2_X1 U430 ( .A(n348), .B(a[2]), .Z(n219) );
  XNOR2_X1 U431 ( .A(n347), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U432 ( .A(n285), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U433 ( .A(n286), .B(n347), .ZN(n198) );
  NAND2_X1 U434 ( .A1(n28), .A2(n342), .ZN(n21) );
  NOR2_X1 U435 ( .A1(n35), .A2(n324), .ZN(n28) );
  INV_X1 U436 ( .A(n322), .ZN(n73) );
  AOI21_X1 U437 ( .B1(n29), .B2(n342), .A(n24), .ZN(n22) );
  AOI21_X1 U438 ( .B1(n37), .B2(n321), .A(n29), .ZN(n27) );
  OAI21_X1 U439 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  XNOR2_X1 U440 ( .A(n8), .B(n55), .ZN(product[5]) );
  INV_X1 U441 ( .A(n303), .ZN(n46) );
  XNOR2_X1 U442 ( .A(n285), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U443 ( .A(n284), .B(b[3]), .ZN(n177) );
  INV_X1 U444 ( .A(n340), .ZN(n75) );
  OAI22_X1 U445 ( .A1(n173), .A2(n283), .B1(n173), .B2(n349), .ZN(n125) );
  OAI22_X1 U446 ( .A1(n283), .A2(n174), .B1(n173), .B2(n349), .ZN(n83) );
  NOR2_X1 U447 ( .A1(n44), .A2(n340), .ZN(n39) );
  OAI21_X1 U448 ( .B1(n45), .B2(n41), .A(n42), .ZN(n40) );
  NAND2_X1 U449 ( .A1(n102), .A2(n107), .ZN(n42) );
  OAI22_X1 U450 ( .A1(n283), .A2(n175), .B1(n174), .B2(n349), .ZN(n142) );
  OAI22_X1 U451 ( .A1(n283), .A2(n176), .B1(n175), .B2(n349), .ZN(n143) );
  OAI22_X1 U452 ( .A1(n283), .A2(n177), .B1(n176), .B2(n349), .ZN(n144) );
  XNOR2_X1 U453 ( .A(n304), .B(b[7]), .ZN(n182) );
  OAI22_X1 U454 ( .A1(n283), .A2(n179), .B1(n178), .B2(n349), .ZN(n146) );
  OAI22_X1 U455 ( .A1(n283), .A2(n178), .B1(n177), .B2(n349), .ZN(n145) );
  XNOR2_X1 U456 ( .A(n291), .B(b[2]), .ZN(n187) );
  OAI22_X1 U457 ( .A1(n221), .A2(n229), .B1(n181), .B2(n225), .ZN(n137) );
  XNOR2_X1 U458 ( .A(n291), .B(b[5]), .ZN(n184) );
  OAI22_X1 U459 ( .A1(n221), .A2(n180), .B1(n179), .B2(n225), .ZN(n147) );
  XNOR2_X1 U460 ( .A(n286), .B(n304), .ZN(n189) );
  XNOR2_X1 U461 ( .A(n304), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U462 ( .A(n291), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U463 ( .A(n291), .B(b[4]), .ZN(n185) );
  INV_X1 U464 ( .A(n234), .ZN(n230) );
  XOR2_X1 U465 ( .A(n7), .B(n274), .Z(product[6]) );
  INV_X1 U466 ( .A(n15), .ZN(n70) );
  OAI21_X1 U467 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  XNOR2_X1 U468 ( .A(n304), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U469 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U470 ( .A(n285), .B(b[1]), .ZN(n197) );
  OAI22_X1 U471 ( .A1(n182), .A2(n287), .B1(n182), .B2(n292), .ZN(n128) );
  OAI22_X1 U472 ( .A1(n287), .A2(n188), .B1(n187), .B2(n292), .ZN(n154) );
  OAI22_X1 U473 ( .A1(n287), .A2(n183), .B1(n182), .B2(n292), .ZN(n89) );
  OAI22_X1 U474 ( .A1(n334), .A2(n187), .B1(n186), .B2(n292), .ZN(n153) );
  OAI22_X1 U475 ( .A1(n287), .A2(n185), .B1(n184), .B2(n292), .ZN(n151) );
  OAI22_X1 U476 ( .A1(n287), .A2(n186), .B1(n185), .B2(n292), .ZN(n152) );
  OAI22_X1 U477 ( .A1(n222), .A2(n184), .B1(n183), .B2(n292), .ZN(n150) );
  INV_X1 U478 ( .A(n292), .ZN(n129) );
  OAI22_X1 U479 ( .A1(n222), .A2(n230), .B1(n190), .B2(n292), .ZN(n138) );
  OAI22_X1 U480 ( .A1(n222), .A2(n189), .B1(n188), .B2(n292), .ZN(n155) );
  OAI21_X1 U481 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U482 ( .B1(n39), .B2(n47), .A(n40), .ZN(n38) );
  XNOR2_X1 U483 ( .A(n20), .B(n1), .ZN(product[12]) );
  INV_X1 U484 ( .A(n338), .ZN(n37) );
  AOI21_X1 U485 ( .B1(n20), .B2(n344), .A(n17), .ZN(n15) );
  OAI22_X1 U486 ( .A1(n326), .A2(n193), .B1(n192), .B2(n296), .ZN(n158) );
  OAI22_X1 U487 ( .A1(n325), .A2(n195), .B1(n194), .B2(n296), .ZN(n160) );
  OAI22_X1 U488 ( .A1(n326), .A2(n194), .B1(n350), .B2(n193), .ZN(n159) );
  OAI22_X1 U489 ( .A1(n325), .A2(n196), .B1(n195), .B2(n296), .ZN(n161) );
  OAI22_X1 U490 ( .A1(n325), .A2(n231), .B1(n199), .B2(n296), .ZN(n139) );
  OAI22_X1 U491 ( .A1(n325), .A2(n197), .B1(n196), .B2(n296), .ZN(n162) );
  OAI22_X1 U492 ( .A1(n326), .A2(n192), .B1(n191), .B2(n296), .ZN(n99) );
  OAI22_X1 U493 ( .A1(n191), .A2(n223), .B1(n191), .B2(n296), .ZN(n131) );
  XNOR2_X1 U494 ( .A(n294), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U495 ( .A(n294), .B(b[6]), .ZN(n201) );
  INV_X1 U496 ( .A(n350), .ZN(n132) );
  OAI22_X1 U497 ( .A1(n223), .A2(n198), .B1(n197), .B2(n350), .ZN(n163) );
  XNOR2_X1 U498 ( .A(n293), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U499 ( .A(n293), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U500 ( .A(n286), .B(n294), .ZN(n207) );
  XNOR2_X1 U501 ( .A(n293), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U502 ( .A(n294), .B(b[3]), .ZN(n204) );
  XNOR2_X1 U503 ( .A(n293), .B(b[1]), .ZN(n206) );
  INV_X1 U504 ( .A(n294), .ZN(n232) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n31, n32, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n73,
         n74, n76, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n128,
         n129, n131, n132, n134, n135, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n216, n217, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n229, n230, n231, n232, n233, n234, n235, n236, n244, n274, n275,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n329, n330, n331, n332,
         n333, n334, n335;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U101 ( .A(n150), .B(n321), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n145), .B(n151), .CI(n100), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n166), .B(n159), .CI(n153), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  BUF_X2 U237 ( .A(n235), .Z(n290) );
  XNOR2_X1 U238 ( .A(n158), .B(n146), .ZN(n106) );
  OR2_X1 U239 ( .A1(n172), .A2(n140), .ZN(n274) );
  NAND3_X1 U240 ( .A1(n70), .A2(n85), .A3(n83), .ZN(n275) );
  BUF_X2 U241 ( .A(n234), .Z(n329) );
  AND3_X1 U242 ( .A1(n275), .A2(n317), .A3(n316), .ZN(product[15]) );
  CLKBUF_X1 U243 ( .A(n45), .Z(n277) );
  XOR2_X1 U244 ( .A(n330), .B(a[4]), .Z(n278) );
  XNOR2_X1 U245 ( .A(n279), .B(n94), .ZN(n92) );
  XNOR2_X1 U246 ( .A(n97), .B(n144), .ZN(n279) );
  CLKBUF_X1 U247 ( .A(n225), .Z(n334) );
  CLKBUF_X1 U248 ( .A(n216), .Z(n292) );
  CLKBUF_X1 U249 ( .A(n216), .Z(n335) );
  AOI21_X1 U250 ( .B1(n327), .B2(n55), .A(n52), .ZN(n280) );
  CLKBUF_X1 U251 ( .A(n44), .Z(n281) );
  INV_X1 U252 ( .A(n34), .ZN(n282) );
  XNOR2_X1 U253 ( .A(n104), .B(n295), .ZN(n283) );
  CLKBUF_X1 U254 ( .A(n330), .Z(n284) );
  OR2_X1 U255 ( .A1(n114), .A2(n117), .ZN(n285) );
  NAND2_X1 U256 ( .A1(n278), .A2(n226), .ZN(n286) );
  OAI21_X1 U257 ( .B1(n299), .B2(n282), .A(n31), .ZN(n287) );
  XOR2_X1 U258 ( .A(n233), .B(a[6]), .Z(n288) );
  XOR2_X1 U259 ( .A(n233), .B(a[6]), .Z(n289) );
  OAI21_X1 U260 ( .B1(n306), .B2(n277), .A(n42), .ZN(n291) );
  NAND2_X1 U261 ( .A1(n96), .A2(n101), .ZN(n36) );
  AOI21_X1 U262 ( .B1(n327), .B2(n55), .A(n52), .ZN(n50) );
  NAND2_X1 U263 ( .A1(n108), .A2(n113), .ZN(n45) );
  NAND2_X1 U264 ( .A1(n220), .A2(n244), .ZN(n293) );
  BUF_X2 U265 ( .A(n236), .Z(n294) );
  NAND2_X1 U266 ( .A1(n220), .A2(n244), .ZN(n224) );
  XNOR2_X1 U267 ( .A(n104), .B(n295), .ZN(n102) );
  XNOR2_X1 U268 ( .A(n109), .B(n106), .ZN(n295) );
  NAND2_X1 U269 ( .A1(n94), .A2(n97), .ZN(n296) );
  NAND2_X1 U270 ( .A1(n94), .A2(n144), .ZN(n297) );
  NAND2_X1 U271 ( .A1(n97), .A2(n144), .ZN(n298) );
  NAND3_X1 U272 ( .A1(n296), .A2(n297), .A3(n298), .ZN(n91) );
  OR2_X1 U273 ( .A1(n88), .A2(n91), .ZN(n324) );
  NOR2_X1 U274 ( .A1(n92), .A2(n95), .ZN(n299) );
  NOR2_X1 U275 ( .A1(n92), .A2(n95), .ZN(n300) );
  NOR2_X1 U276 ( .A1(n35), .A2(n300), .ZN(n301) );
  NAND2_X1 U277 ( .A1(n104), .A2(n109), .ZN(n302) );
  NAND2_X1 U278 ( .A1(n104), .A2(n106), .ZN(n303) );
  NAND2_X1 U279 ( .A1(n109), .A2(n106), .ZN(n304) );
  NAND3_X1 U280 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n101) );
  XNOR2_X1 U281 ( .A(n232), .B(n135), .ZN(n220) );
  XNOR2_X1 U282 ( .A(n329), .B(a[6]), .ZN(n305) );
  NOR2_X1 U283 ( .A1(n102), .A2(n107), .ZN(n306) );
  NAND2_X1 U284 ( .A1(n217), .A2(n305), .ZN(n307) );
  NAND2_X1 U285 ( .A1(n289), .A2(n305), .ZN(n308) );
  NAND2_X1 U286 ( .A1(n288), .A2(n305), .ZN(n221) );
  CLKBUF_X1 U287 ( .A(n70), .Z(n309) );
  NAND3_X1 U288 ( .A1(n312), .A2(n314), .A3(n313), .ZN(n310) );
  XOR2_X1 U289 ( .A(n85), .B(n84), .Z(n311) );
  XOR2_X1 U290 ( .A(n311), .B(n309), .Z(product[13]) );
  NAND2_X1 U291 ( .A1(n85), .A2(n84), .ZN(n312) );
  NAND2_X1 U292 ( .A1(n85), .A2(n70), .ZN(n313) );
  NAND2_X1 U293 ( .A1(n70), .A2(n84), .ZN(n314) );
  NAND3_X1 U294 ( .A1(n312), .A2(n313), .A3(n314), .ZN(n14) );
  XOR2_X1 U295 ( .A(n141), .B(n83), .Z(n315) );
  XOR2_X1 U296 ( .A(n315), .B(n310), .Z(product[14]) );
  NAND2_X1 U297 ( .A1(n141), .A2(n83), .ZN(n316) );
  NAND2_X1 U298 ( .A1(n14), .A2(n141), .ZN(n317) );
  NAND2_X1 U299 ( .A1(n278), .A2(n226), .ZN(n318) );
  NAND2_X1 U300 ( .A1(n323), .A2(n226), .ZN(n222) );
  OAI21_X1 U301 ( .B1(n48), .B2(n280), .A(n49), .ZN(n319) );
  CLKBUF_X1 U302 ( .A(n20), .Z(n320) );
  OAI22_X1 U303 ( .A1(n223), .A2(n192), .B1(n191), .B2(n332), .ZN(n321) );
  AOI21_X1 U304 ( .B1(n39), .B2(n319), .A(n291), .ZN(n322) );
  NOR2_X1 U305 ( .A1(n108), .A2(n113), .ZN(n44) );
  INV_X2 U306 ( .A(n135), .ZN(n244) );
  XOR2_X1 U307 ( .A(n329), .B(a[4]), .Z(n323) );
  XNOR2_X1 U308 ( .A(n37), .B(n4), .ZN(product[9]) );
  INV_X1 U309 ( .A(n35), .ZN(n74) );
  INV_X1 U310 ( .A(n26), .ZN(n24) );
  NAND2_X1 U311 ( .A1(n326), .A2(n19), .ZN(n1) );
  XOR2_X1 U312 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U313 ( .A1(n73), .A2(n31), .ZN(n3) );
  AOI21_X1 U314 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  INV_X1 U315 ( .A(n300), .ZN(n73) );
  XOR2_X1 U316 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U317 ( .A1(n76), .A2(n277), .ZN(n6) );
  INV_X1 U318 ( .A(n281), .ZN(n76) );
  XOR2_X1 U319 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U320 ( .A1(n324), .A2(n26), .ZN(n2) );
  XNOR2_X1 U321 ( .A(n8), .B(n55), .ZN(product[5]) );
  XNOR2_X1 U322 ( .A(n43), .B(n5), .ZN(product[8]) );
  OAI21_X1 U323 ( .B1(n46), .B2(n281), .A(n277), .ZN(n43) );
  XNOR2_X1 U324 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U325 ( .A1(n325), .A2(n66), .ZN(n11) );
  NAND2_X1 U326 ( .A1(n285), .A2(n49), .ZN(n7) );
  INV_X1 U327 ( .A(n19), .ZN(n17) );
  XOR2_X1 U328 ( .A(n10), .B(n62), .Z(product[3]) );
  NAND2_X1 U329 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U330 ( .A(n60), .ZN(n80) );
  XOR2_X1 U331 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U332 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U333 ( .A(n56), .ZN(n79) );
  OR2_X1 U334 ( .A1(n158), .A2(n146), .ZN(n105) );
  NOR2_X1 U335 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U336 ( .A(n83), .ZN(n84) );
  NAND2_X1 U337 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U338 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U339 ( .A1(n114), .A2(n117), .ZN(n49) );
  OR2_X1 U340 ( .A1(n171), .A2(n164), .ZN(n325) );
  NAND2_X1 U341 ( .A1(n92), .A2(n95), .ZN(n31) );
  OR2_X1 U342 ( .A1(n87), .A2(n86), .ZN(n326) );
  OR2_X1 U343 ( .A1(n118), .A2(n121), .ZN(n327) );
  AND2_X1 U344 ( .A1(n335), .A2(n132), .ZN(n164) );
  AND2_X1 U345 ( .A1(n292), .A2(n126), .ZN(n148) );
  INV_X1 U346 ( .A(n128), .ZN(n149) );
  INV_X1 U347 ( .A(n89), .ZN(n90) );
  AND2_X1 U348 ( .A1(n292), .A2(n129), .ZN(n156) );
  OAI22_X1 U349 ( .A1(n293), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OR2_X1 U350 ( .A1(n216), .A2(n230), .ZN(n190) );
  BUF_X2 U351 ( .A(n226), .Z(n331) );
  OAI22_X1 U352 ( .A1(n293), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  NOR2_X1 U353 ( .A1(n122), .A2(n123), .ZN(n56) );
  INV_X1 U354 ( .A(n125), .ZN(n141) );
  NAND2_X1 U355 ( .A1(n122), .A2(n123), .ZN(n57) );
  INV_X1 U356 ( .A(n99), .ZN(n100) );
  OR2_X1 U357 ( .A1(n335), .A2(n229), .ZN(n181) );
  AND2_X1 U358 ( .A1(n274), .A2(n69), .ZN(product[1]) );
  OR2_X1 U359 ( .A1(n335), .A2(n231), .ZN(n199) );
  OAI22_X1 U360 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI22_X1 U361 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U362 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  OR2_X1 U363 ( .A1(n292), .A2(n232), .ZN(n208) );
  AND2_X1 U364 ( .A1(n216), .A2(n135), .ZN(product[0]) );
  NAND2_X1 U365 ( .A1(n171), .A2(n164), .ZN(n66) );
  CLKBUF_X3 U366 ( .A(n234), .Z(n330) );
  XNOR2_X1 U367 ( .A(n235), .B(a[4]), .ZN(n226) );
  BUF_X2 U368 ( .A(n227), .Z(n332) );
  XNOR2_X1 U369 ( .A(n236), .B(a[2]), .ZN(n227) );
  INV_X1 U370 ( .A(n233), .ZN(n229) );
  XNOR2_X1 U371 ( .A(n292), .B(n233), .ZN(n180) );
  XNOR2_X1 U372 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U373 ( .A(n233), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U374 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U375 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U376 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U377 ( .A(n233), .B(b[7]), .ZN(n173) );
  NOR2_X1 U378 ( .A1(n124), .A2(n139), .ZN(n60) );
  OAI22_X1 U379 ( .A1(n293), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U380 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  NAND2_X1 U381 ( .A1(n74), .A2(n282), .ZN(n4) );
  INV_X1 U382 ( .A(n36), .ZN(n34) );
  NAND2_X1 U383 ( .A1(n327), .A2(n54), .ZN(n8) );
  NAND2_X1 U384 ( .A1(n333), .A2(n42), .ZN(n5) );
  INV_X1 U385 ( .A(n134), .ZN(n165) );
  OAI22_X1 U386 ( .A1(n200), .A2(n293), .B1(n200), .B2(n244), .ZN(n134) );
  OR2_X1 U387 ( .A1(n283), .A2(n107), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n329), .B(a[6]), .ZN(n225) );
  NOR2_X1 U389 ( .A1(n102), .A2(n107), .ZN(n41) );
  XOR2_X1 U390 ( .A(n233), .B(a[6]), .Z(n217) );
  OAI21_X1 U391 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  AOI21_X1 U392 ( .B1(n325), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U393 ( .A(n69), .ZN(n67) );
  INV_X1 U394 ( .A(n66), .ZN(n64) );
  OAI22_X1 U395 ( .A1(n293), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  NAND2_X1 U396 ( .A1(n118), .A2(n121), .ZN(n54) );
  NAND2_X1 U397 ( .A1(n28), .A2(n324), .ZN(n21) );
  INV_X1 U398 ( .A(n131), .ZN(n157) );
  NAND2_X1 U399 ( .A1(n283), .A2(n107), .ZN(n42) );
  INV_X1 U400 ( .A(n54), .ZN(n52) );
  INV_X1 U401 ( .A(n59), .ZN(n58) );
  OAI21_X1 U402 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  AOI21_X1 U403 ( .B1(n29), .B2(n324), .A(n24), .ZN(n22) );
  AOI21_X1 U404 ( .B1(n37), .B2(n301), .A(n287), .ZN(n27) );
  OAI21_X1 U405 ( .B1(n299), .B2(n36), .A(n31), .ZN(n29) );
  NOR2_X1 U406 ( .A1(n35), .A2(n300), .ZN(n28) );
  NOR2_X1 U407 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U408 ( .A1(n124), .A2(n139), .ZN(n61) );
  OAI21_X1 U409 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  OAI21_X1 U410 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  INV_X1 U411 ( .A(n319), .ZN(n46) );
  AOI21_X1 U412 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U413 ( .A1(n172), .A2(n140), .ZN(n69) );
  XNOR2_X1 U414 ( .A(n294), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U415 ( .A(n294), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U416 ( .A(n294), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U417 ( .A(n294), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U418 ( .A(n294), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U419 ( .A(n294), .B(b[3]), .ZN(n204) );
  XNOR2_X1 U420 ( .A(n216), .B(n294), .ZN(n207) );
  INV_X1 U421 ( .A(n236), .ZN(n232) );
  XOR2_X1 U422 ( .A(n7), .B(n280), .Z(product[6]) );
  OAI22_X1 U423 ( .A1(n182), .A2(n286), .B1(n182), .B2(n331), .ZN(n128) );
  OAI22_X1 U424 ( .A1(n286), .A2(n188), .B1(n187), .B2(n331), .ZN(n154) );
  OAI22_X1 U425 ( .A1(n286), .A2(n183), .B1(n182), .B2(n331), .ZN(n89) );
  OAI22_X1 U426 ( .A1(n286), .A2(n186), .B1(n185), .B2(n331), .ZN(n152) );
  OAI22_X1 U427 ( .A1(n318), .A2(n187), .B1(n186), .B2(n331), .ZN(n153) );
  OAI22_X1 U428 ( .A1(n318), .A2(n185), .B1(n184), .B2(n331), .ZN(n151) );
  OAI22_X1 U429 ( .A1(n286), .A2(n184), .B1(n183), .B2(n331), .ZN(n150) );
  INV_X1 U430 ( .A(n331), .ZN(n129) );
  XNOR2_X1 U431 ( .A(n290), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U432 ( .A(n290), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U433 ( .A(n290), .B(b[3]), .ZN(n195) );
  OAI22_X1 U434 ( .A1(n222), .A2(n230), .B1(n190), .B2(n331), .ZN(n138) );
  OAI22_X1 U435 ( .A1(n222), .A2(n189), .B1(n188), .B2(n331), .ZN(n155) );
  XNOR2_X1 U436 ( .A(n290), .B(b[2]), .ZN(n196) );
  INV_X1 U437 ( .A(n290), .ZN(n231) );
  XNOR2_X1 U438 ( .A(n290), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U439 ( .A(n290), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U440 ( .A(n335), .B(n290), .ZN(n198) );
  XOR2_X1 U441 ( .A(n235), .B(a[2]), .Z(n219) );
  INV_X1 U442 ( .A(n15), .ZN(n70) );
  OAI22_X1 U443 ( .A1(n173), .A2(n307), .B1(n173), .B2(n334), .ZN(n125) );
  OAI22_X1 U444 ( .A1(n308), .A2(n174), .B1(n173), .B2(n334), .ZN(n83) );
  NOR2_X1 U445 ( .A1(n306), .A2(n44), .ZN(n39) );
  OAI21_X1 U446 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI22_X1 U447 ( .A1(n307), .A2(n175), .B1(n174), .B2(n334), .ZN(n142) );
  OAI22_X1 U448 ( .A1(n308), .A2(n176), .B1(n175), .B2(n334), .ZN(n143) );
  OAI22_X1 U449 ( .A1(n307), .A2(n177), .B1(n176), .B2(n334), .ZN(n144) );
  XNOR2_X1 U450 ( .A(n284), .B(b[7]), .ZN(n182) );
  OAI22_X1 U451 ( .A1(n307), .A2(n178), .B1(n177), .B2(n225), .ZN(n145) );
  INV_X1 U452 ( .A(n225), .ZN(n126) );
  OAI22_X1 U453 ( .A1(n308), .A2(n179), .B1(n178), .B2(n225), .ZN(n146) );
  XNOR2_X1 U454 ( .A(n330), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U455 ( .A(n330), .B(b[5]), .ZN(n184) );
  OAI22_X1 U456 ( .A1(n221), .A2(n229), .B1(n181), .B2(n225), .ZN(n137) );
  OAI22_X1 U457 ( .A1(n221), .A2(n180), .B1(n179), .B2(n225), .ZN(n147) );
  XNOR2_X1 U458 ( .A(n284), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U459 ( .A(n330), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U460 ( .A(n330), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U461 ( .A(n335), .B(n330), .ZN(n189) );
  INV_X1 U462 ( .A(n330), .ZN(n230) );
  XNOR2_X1 U463 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U464 ( .A(n330), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U465 ( .A(n290), .B(b[1]), .ZN(n197) );
  XNOR2_X1 U466 ( .A(n294), .B(b[1]), .ZN(n206) );
  XNOR2_X1 U467 ( .A(n320), .B(n1), .ZN(product[12]) );
  INV_X1 U468 ( .A(n322), .ZN(n37) );
  AOI21_X1 U469 ( .B1(n20), .B2(n326), .A(n17), .ZN(n15) );
  OAI22_X1 U470 ( .A1(n223), .A2(n193), .B1(n192), .B2(n332), .ZN(n158) );
  OAI22_X1 U471 ( .A1(n223), .A2(n195), .B1(n194), .B2(n332), .ZN(n160) );
  OAI22_X1 U472 ( .A1(n223), .A2(n194), .B1(n193), .B2(n332), .ZN(n159) );
  OAI22_X1 U473 ( .A1(n223), .A2(n196), .B1(n195), .B2(n332), .ZN(n161) );
  OAI22_X1 U474 ( .A1(n223), .A2(n231), .B1(n199), .B2(n332), .ZN(n139) );
  OAI22_X1 U475 ( .A1(n223), .A2(n197), .B1(n196), .B2(n332), .ZN(n162) );
  OAI22_X1 U476 ( .A1(n223), .A2(n192), .B1(n191), .B2(n332), .ZN(n99) );
  OAI22_X1 U477 ( .A1(n191), .A2(n223), .B1(n191), .B2(n332), .ZN(n131) );
  INV_X1 U478 ( .A(n332), .ZN(n132) );
  OAI22_X1 U479 ( .A1(n223), .A2(n198), .B1(n197), .B2(n332), .ZN(n163) );
  NAND2_X2 U480 ( .A1(n219), .A2(n227), .ZN(n223) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70,
         n74, n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n128, n129, n131, n132, n134, n135, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n216, n217, n218, n220, n221, n222, n223, n224, n225,
         n226, n229, n230, n231, n232, n233, n234, n235, n236, n244, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342,
         n343, n344;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n157), .B(n295), .CI(n150), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n100), .B(n145), .CI(n151), .CO(n97), .S(n98) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n159), .B(n166), .CI(n153), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n137), .B(n147), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  BUF_X2 U237 ( .A(n216), .Z(n344) );
  BUF_X1 U238 ( .A(n235), .Z(n274) );
  OR2_X1 U239 ( .A1(n172), .A2(n140), .ZN(n275) );
  NAND2_X1 U240 ( .A1(n338), .A2(n218), .ZN(n276) );
  CLKBUF_X1 U241 ( .A(n236), .Z(n277) );
  INV_X1 U242 ( .A(n230), .ZN(n278) );
  BUF_X2 U243 ( .A(n340), .Z(n287) );
  INV_X1 U244 ( .A(n34), .ZN(n279) );
  NOR2_X1 U245 ( .A1(n30), .A2(n35), .ZN(n280) );
  CLKBUF_X1 U246 ( .A(n44), .Z(n281) );
  CLKBUF_X1 U247 ( .A(n47), .Z(n282) );
  OR2_X2 U248 ( .A1(n327), .A2(n328), .ZN(n223) );
  OAI22_X1 U249 ( .A1(n290), .A2(n186), .B1(n185), .B2(n339), .ZN(n283) );
  AND3_X1 U250 ( .A1(n70), .A2(n85), .A3(n83), .ZN(n284) );
  INV_X1 U251 ( .A(n284), .ZN(n315) );
  CLKBUF_X1 U252 ( .A(n92), .Z(n285) );
  BUF_X2 U253 ( .A(n340), .Z(n286) );
  XOR2_X1 U254 ( .A(n233), .B(a[6]), .Z(n288) );
  OR2_X2 U255 ( .A1(n327), .A2(n328), .ZN(n289) );
  NAND2_X1 U256 ( .A1(n338), .A2(n218), .ZN(n290) );
  NAND2_X1 U257 ( .A1(n338), .A2(n218), .ZN(n341) );
  CLKBUF_X1 U258 ( .A(n236), .Z(n291) );
  CLKBUF_X1 U259 ( .A(n45), .Z(n292) );
  XNOR2_X2 U260 ( .A(n234), .B(a[6]), .ZN(n225) );
  AOI21_X1 U261 ( .B1(n333), .B2(n55), .A(n52), .ZN(n50) );
  CLKBUF_X1 U262 ( .A(n343), .Z(n293) );
  NOR2_X1 U263 ( .A1(n92), .A2(n95), .ZN(n294) );
  OAI22_X1 U264 ( .A1(n289), .A2(n192), .B1(n191), .B2(n287), .ZN(n295) );
  CLKBUF_X1 U265 ( .A(n35), .Z(n296) );
  XNOR2_X1 U266 ( .A(n297), .B(n111), .ZN(n104) );
  XNOR2_X1 U267 ( .A(n165), .B(n152), .ZN(n297) );
  CLKBUF_X1 U268 ( .A(n70), .Z(n298) );
  OAI21_X1 U269 ( .B1(n41), .B2(n45), .A(n42), .ZN(n299) );
  NAND3_X1 U270 ( .A1(n311), .A2(n310), .A3(n312), .ZN(n300) );
  CLKBUF_X1 U271 ( .A(n29), .Z(n301) );
  XOR2_X1 U272 ( .A(n168), .B(n161), .Z(n302) );
  XOR2_X1 U273 ( .A(n120), .B(n302), .Z(n118) );
  NAND2_X1 U274 ( .A1(n120), .A2(n168), .ZN(n303) );
  NAND2_X1 U275 ( .A1(n120), .A2(n161), .ZN(n304) );
  NAND2_X1 U276 ( .A1(n168), .A2(n161), .ZN(n305) );
  NAND3_X1 U277 ( .A1(n303), .A2(n304), .A3(n305), .ZN(n117) );
  XNOR2_X1 U278 ( .A(n306), .B(n300), .ZN(product[14]) );
  XNOR2_X1 U279 ( .A(n141), .B(n83), .ZN(n306) );
  AND3_X1 U280 ( .A1(n314), .A2(n315), .A3(n313), .ZN(product[15]) );
  BUF_X2 U281 ( .A(n226), .Z(n338) );
  NAND2_X1 U282 ( .A1(n108), .A2(n113), .ZN(n45) );
  XNOR2_X1 U283 ( .A(n104), .B(n308), .ZN(n102) );
  XNOR2_X1 U284 ( .A(n109), .B(n106), .ZN(n308) );
  XOR2_X1 U285 ( .A(n85), .B(n84), .Z(n309) );
  XOR2_X1 U286 ( .A(n309), .B(n298), .Z(product[13]) );
  NAND2_X1 U287 ( .A1(n85), .A2(n84), .ZN(n310) );
  NAND2_X1 U288 ( .A1(n70), .A2(n85), .ZN(n311) );
  NAND2_X1 U289 ( .A1(n70), .A2(n84), .ZN(n312) );
  NAND3_X1 U290 ( .A1(n312), .A2(n311), .A3(n310), .ZN(n14) );
  NAND2_X1 U291 ( .A1(n141), .A2(n83), .ZN(n313) );
  NAND2_X1 U292 ( .A1(n14), .A2(n141), .ZN(n314) );
  NAND2_X1 U293 ( .A1(n165), .A2(n283), .ZN(n316) );
  NAND2_X1 U294 ( .A1(n165), .A2(n111), .ZN(n317) );
  NAND2_X1 U295 ( .A1(n283), .A2(n111), .ZN(n318) );
  NAND3_X1 U296 ( .A1(n316), .A2(n317), .A3(n318), .ZN(n103) );
  NAND2_X1 U297 ( .A1(n109), .A2(n106), .ZN(n319) );
  NAND2_X1 U298 ( .A1(n109), .A2(n104), .ZN(n320) );
  NAND2_X1 U299 ( .A1(n106), .A2(n104), .ZN(n321) );
  NAND3_X1 U300 ( .A1(n319), .A2(n320), .A3(n321), .ZN(n101) );
  CLKBUF_X2 U301 ( .A(n226), .Z(n339) );
  NAND2_X1 U302 ( .A1(n236), .A2(n322), .ZN(n323) );
  NAND2_X1 U303 ( .A1(n232), .A2(n135), .ZN(n324) );
  NAND2_X1 U304 ( .A1(n323), .A2(n324), .ZN(n220) );
  INV_X1 U305 ( .A(n135), .ZN(n322) );
  NAND2_X2 U306 ( .A1(n220), .A2(n244), .ZN(n325) );
  NAND2_X1 U307 ( .A1(n220), .A2(n244), .ZN(n224) );
  OR2_X1 U308 ( .A1(n285), .A2(n95), .ZN(n326) );
  XNOR2_X1 U309 ( .A(n235), .B(a[2]), .ZN(n327) );
  XOR2_X1 U310 ( .A(n236), .B(a[2]), .Z(n328) );
  CLKBUF_X1 U311 ( .A(n20), .Z(n329) );
  AOI21_X1 U312 ( .B1(n39), .B2(n282), .A(n299), .ZN(n330) );
  XNOR2_X1 U313 ( .A(n234), .B(a[6]), .ZN(n331) );
  NOR2_X1 U314 ( .A1(n102), .A2(n107), .ZN(n332) );
  INV_X1 U315 ( .A(n296), .ZN(n74) );
  XNOR2_X1 U316 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U317 ( .A1(n74), .A2(n279), .ZN(n4) );
  INV_X1 U318 ( .A(n36), .ZN(n34) );
  INV_X1 U319 ( .A(n54), .ZN(n52) );
  INV_X1 U320 ( .A(n26), .ZN(n24) );
  OAI21_X1 U321 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  INV_X1 U322 ( .A(n59), .ZN(n58) );
  NOR2_X1 U323 ( .A1(n102), .A2(n107), .ZN(n41) );
  NAND2_X1 U324 ( .A1(n336), .A2(n19), .ZN(n1) );
  XOR2_X1 U325 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U326 ( .A1(n326), .A2(n31), .ZN(n3) );
  AOI21_X1 U327 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U328 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U329 ( .A1(n76), .A2(n292), .ZN(n6) );
  INV_X1 U330 ( .A(n281), .ZN(n76) );
  XOR2_X1 U331 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U332 ( .A1(n335), .A2(n26), .ZN(n2) );
  NAND2_X1 U333 ( .A1(n102), .A2(n107), .ZN(n42) );
  XNOR2_X1 U334 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U335 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U336 ( .B1(n46), .B2(n281), .A(n292), .ZN(n43) );
  XNOR2_X1 U337 ( .A(n8), .B(n55), .ZN(product[5]) );
  NAND2_X1 U338 ( .A1(n333), .A2(n54), .ZN(n8) );
  XNOR2_X1 U339 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U340 ( .A1(n334), .A2(n66), .ZN(n11) );
  NAND2_X1 U341 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U342 ( .A(n48), .ZN(n77) );
  NAND2_X1 U343 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U344 ( .A(n60), .ZN(n80) );
  XOR2_X1 U345 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U346 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U347 ( .A(n56), .ZN(n79) );
  INV_X1 U348 ( .A(n19), .ZN(n17) );
  NOR2_X1 U349 ( .A1(n108), .A2(n113), .ZN(n44) );
  XNOR2_X1 U350 ( .A(n158), .B(n146), .ZN(n106) );
  NOR2_X1 U351 ( .A1(n92), .A2(n95), .ZN(n30) );
  OR2_X1 U352 ( .A1(n118), .A2(n121), .ZN(n333) );
  OR2_X1 U353 ( .A1(n171), .A2(n164), .ZN(n334) );
  NOR2_X1 U354 ( .A1(n122), .A2(n123), .ZN(n56) );
  OR2_X1 U355 ( .A1(n158), .A2(n146), .ZN(n105) );
  NOR2_X1 U356 ( .A1(n114), .A2(n117), .ZN(n48) );
  NOR2_X1 U357 ( .A1(n124), .A2(n139), .ZN(n60) );
  INV_X1 U358 ( .A(n83), .ZN(n84) );
  OR2_X1 U359 ( .A1(n88), .A2(n91), .ZN(n335) );
  NAND2_X1 U360 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U361 ( .A1(n87), .A2(n86), .ZN(n19) );
  INV_X1 U362 ( .A(n69), .ZN(n67) );
  NAND2_X1 U363 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U364 ( .A1(n122), .A2(n123), .ZN(n57) );
  OR2_X1 U365 ( .A1(n87), .A2(n86), .ZN(n336) );
  OR2_X1 U366 ( .A1(n344), .A2(n231), .ZN(n199) );
  INV_X1 U367 ( .A(n128), .ZN(n149) );
  INV_X1 U368 ( .A(n89), .ZN(n90) );
  AND2_X1 U369 ( .A1(n344), .A2(n129), .ZN(n156) );
  AND2_X1 U370 ( .A1(n344), .A2(n126), .ZN(n148) );
  INV_X1 U371 ( .A(n125), .ZN(n141) );
  OR2_X1 U372 ( .A1(n344), .A2(n229), .ZN(n181) );
  AND2_X1 U373 ( .A1(n275), .A2(n69), .ZN(product[1]) );
  INV_X1 U374 ( .A(n134), .ZN(n165) );
  AND2_X1 U375 ( .A1(n344), .A2(n132), .ZN(n164) );
  OR2_X1 U376 ( .A1(n344), .A2(n230), .ZN(n190) );
  XNOR2_X1 U377 ( .A(n236), .B(a[2]), .ZN(n340) );
  OR2_X1 U378 ( .A1(n344), .A2(n232), .ZN(n208) );
  INV_X1 U379 ( .A(n135), .ZN(n244) );
  AND2_X1 U380 ( .A1(n344), .A2(n135), .ZN(product[0]) );
  NAND2_X1 U381 ( .A1(n218), .A2(n338), .ZN(n222) );
  NAND2_X1 U382 ( .A1(n171), .A2(n164), .ZN(n66) );
  XNOR2_X1 U383 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U384 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U385 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U386 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U387 ( .A(n344), .B(n233), .ZN(n180) );
  INV_X1 U388 ( .A(n233), .ZN(n229) );
  XNOR2_X1 U389 ( .A(n235), .B(a[4]), .ZN(n226) );
  XOR2_X1 U390 ( .A(n233), .B(a[6]), .Z(n217) );
  OAI22_X1 U391 ( .A1(n325), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  OAI22_X1 U392 ( .A1(n325), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U393 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U394 ( .A1(n325), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  OAI22_X1 U395 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U396 ( .A1(n325), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI22_X1 U397 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  XOR2_X1 U398 ( .A(n10), .B(n62), .Z(product[3]) );
  OAI21_X1 U399 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  AOI21_X1 U400 ( .B1(n334), .B2(n67), .A(n64), .ZN(n62) );
  NAND2_X1 U401 ( .A1(n172), .A2(n140), .ZN(n69) );
  OAI22_X1 U402 ( .A1(n325), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  NAND2_X1 U403 ( .A1(n28), .A2(n335), .ZN(n21) );
  NOR2_X1 U404 ( .A1(n30), .A2(n35), .ZN(n28) );
  INV_X1 U405 ( .A(n131), .ZN(n157) );
  NAND2_X1 U406 ( .A1(n288), .A2(n331), .ZN(n342) );
  NAND2_X1 U407 ( .A1(n217), .A2(n225), .ZN(n343) );
  NAND2_X1 U408 ( .A1(n217), .A2(n331), .ZN(n221) );
  NOR2_X1 U409 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U410 ( .A1(n96), .A2(n101), .ZN(n36) );
  XNOR2_X1 U411 ( .A(n233), .B(b[3]), .ZN(n177) );
  NAND2_X1 U412 ( .A1(n124), .A2(n139), .ZN(n61) );
  AOI21_X1 U413 ( .B1(n37), .B2(n280), .A(n301), .ZN(n27) );
  AOI21_X1 U414 ( .B1(n29), .B2(n335), .A(n24), .ZN(n22) );
  OAI21_X1 U415 ( .B1(n36), .B2(n294), .A(n31), .ZN(n29) );
  INV_X1 U416 ( .A(n99), .ZN(n100) );
  INV_X1 U417 ( .A(n66), .ZN(n64) );
  OAI22_X1 U418 ( .A1(n325), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  XNOR2_X1 U419 ( .A(n233), .B(b[1]), .ZN(n179) );
  INV_X1 U420 ( .A(n332), .ZN(n75) );
  NOR2_X1 U421 ( .A1(n44), .A2(n332), .ZN(n39) );
  OAI21_X1 U422 ( .B1(n45), .B2(n41), .A(n42), .ZN(n40) );
  XNOR2_X1 U423 ( .A(n233), .B(b[7]), .ZN(n173) );
  NAND2_X1 U424 ( .A1(n92), .A2(n95), .ZN(n31) );
  NAND2_X1 U425 ( .A1(n118), .A2(n121), .ZN(n54) );
  OAI22_X1 U426 ( .A1(n182), .A2(n290), .B1(n182), .B2(n339), .ZN(n128) );
  OAI22_X1 U427 ( .A1(n290), .A2(n188), .B1(n187), .B2(n339), .ZN(n154) );
  OAI22_X1 U428 ( .A1(n290), .A2(n183), .B1(n182), .B2(n339), .ZN(n89) );
  INV_X1 U429 ( .A(n339), .ZN(n129) );
  OAI22_X1 U430 ( .A1(n276), .A2(n187), .B1(n186), .B2(n339), .ZN(n153) );
  OAI22_X1 U431 ( .A1(n290), .A2(n186), .B1(n185), .B2(n339), .ZN(n152) );
  OAI22_X1 U432 ( .A1(n276), .A2(n185), .B1(n184), .B2(n339), .ZN(n151) );
  OAI22_X1 U433 ( .A1(n341), .A2(n184), .B1(n183), .B2(n339), .ZN(n150) );
  OAI22_X1 U434 ( .A1(n222), .A2(n230), .B1(n190), .B2(n339), .ZN(n138) );
  OAI22_X1 U435 ( .A1(n222), .A2(n189), .B1(n188), .B2(n339), .ZN(n155) );
  OAI21_X1 U436 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  XNOR2_X1 U437 ( .A(n278), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U438 ( .A(n234), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U439 ( .A(n234), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U440 ( .A(n234), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U441 ( .A(n344), .B(n234), .ZN(n189) );
  INV_X1 U442 ( .A(n234), .ZN(n230) );
  XNOR2_X1 U443 ( .A(n234), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U444 ( .A(n234), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U445 ( .A(n234), .B(b[1]), .ZN(n188) );
  XOR2_X1 U446 ( .A(n234), .B(a[4]), .Z(n218) );
  XOR2_X1 U447 ( .A(n7), .B(n50), .Z(product[6]) );
  INV_X1 U448 ( .A(n282), .ZN(n46) );
  AOI21_X1 U449 ( .B1(n39), .B2(n47), .A(n40), .ZN(n38) );
  OAI21_X1 U450 ( .B1(n48), .B2(n50), .A(n49), .ZN(n47) );
  XNOR2_X1 U451 ( .A(n274), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U452 ( .A(n274), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U453 ( .A(n274), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U454 ( .A(n274), .B(b[2]), .ZN(n196) );
  INV_X1 U455 ( .A(n274), .ZN(n231) );
  XNOR2_X1 U456 ( .A(n235), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U457 ( .A(n235), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U458 ( .A(n344), .B(n274), .ZN(n198) );
  XNOR2_X1 U459 ( .A(n235), .B(b[1]), .ZN(n197) );
  INV_X1 U460 ( .A(n15), .ZN(n70) );
  OAI22_X1 U461 ( .A1(n173), .A2(n293), .B1(n173), .B2(n225), .ZN(n125) );
  OAI22_X1 U462 ( .A1(n342), .A2(n174), .B1(n173), .B2(n225), .ZN(n83) );
  OAI22_X1 U463 ( .A1(n221), .A2(n175), .B1(n174), .B2(n331), .ZN(n142) );
  OAI22_X1 U464 ( .A1(n342), .A2(n176), .B1(n175), .B2(n225), .ZN(n143) );
  OAI22_X1 U465 ( .A1(n293), .A2(n177), .B1(n176), .B2(n331), .ZN(n144) );
  OAI22_X1 U466 ( .A1(n221), .A2(n179), .B1(n178), .B2(n225), .ZN(n146) );
  OAI22_X1 U467 ( .A1(n343), .A2(n178), .B1(n177), .B2(n225), .ZN(n145) );
  INV_X1 U468 ( .A(n225), .ZN(n126) );
  OAI22_X1 U469 ( .A1(n342), .A2(n229), .B1(n181), .B2(n225), .ZN(n137) );
  OAI22_X1 U470 ( .A1(n221), .A2(n180), .B1(n179), .B2(n225), .ZN(n147) );
  XNOR2_X1 U471 ( .A(n329), .B(n1), .ZN(product[12]) );
  INV_X1 U472 ( .A(n330), .ZN(n37) );
  AOI21_X1 U473 ( .B1(n20), .B2(n336), .A(n17), .ZN(n15) );
  OAI22_X1 U474 ( .A1(n223), .A2(n193), .B1(n192), .B2(n287), .ZN(n158) );
  OAI22_X1 U475 ( .A1(n223), .A2(n195), .B1(n194), .B2(n286), .ZN(n160) );
  OAI22_X1 U476 ( .A1(n223), .A2(n194), .B1(n193), .B2(n286), .ZN(n159) );
  OAI22_X1 U477 ( .A1(n223), .A2(n196), .B1(n195), .B2(n287), .ZN(n161) );
  OAI22_X1 U478 ( .A1(n223), .A2(n231), .B1(n199), .B2(n286), .ZN(n139) );
  OAI22_X1 U479 ( .A1(n223), .A2(n197), .B1(n196), .B2(n286), .ZN(n162) );
  OAI22_X1 U480 ( .A1(n289), .A2(n192), .B1(n191), .B2(n286), .ZN(n99) );
  OAI22_X1 U481 ( .A1(n191), .A2(n289), .B1(n191), .B2(n287), .ZN(n131) );
  XNOR2_X1 U482 ( .A(n291), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U483 ( .A(n277), .B(b[6]), .ZN(n201) );
  INV_X1 U484 ( .A(n286), .ZN(n132) );
  OAI22_X1 U485 ( .A1(n223), .A2(n198), .B1(n197), .B2(n287), .ZN(n163) );
  XNOR2_X1 U486 ( .A(n291), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U487 ( .A(n236), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U488 ( .A(n344), .B(n291), .ZN(n207) );
  XNOR2_X1 U489 ( .A(n277), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U490 ( .A(n277), .B(b[3]), .ZN(n204) );
  XNOR2_X1 U491 ( .A(n277), .B(b[1]), .ZN(n206) );
  INV_X1 U492 ( .A(n236), .ZN(n232) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n73,
         n74, n75, n76, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n129, n131, n132, n134, n135, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n216, n217, n220, n221, n222, n223, n224, n225, n226, n227,
         n229, n230, n231, n232, n233, n234, n235, n236, n244, n274, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U101 ( .A(n150), .B(n312), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n145), .B(n151), .CI(n100), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n153), .B(n166), .CI(n159), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  HA_X1 U115 ( .A(n138), .B(n155), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  BUF_X1 U237 ( .A(n235), .Z(n326) );
  NOR2_X1 U238 ( .A1(n108), .A2(n113), .ZN(n44) );
  OR2_X1 U239 ( .A1(n172), .A2(n140), .ZN(n274) );
  AND3_X1 U240 ( .A1(n281), .A2(n282), .A3(n283), .ZN(product[15]) );
  INV_X1 U241 ( .A(n15), .ZN(n276) );
  CLKBUF_X1 U242 ( .A(n28), .Z(n277) );
  NAND3_X1 U243 ( .A1(n335), .A2(n336), .A3(n337), .ZN(n278) );
  AND3_X1 U244 ( .A1(n276), .A2(n85), .A3(n83), .ZN(n279) );
  INV_X1 U245 ( .A(n279), .ZN(n282) );
  XOR2_X1 U246 ( .A(n141), .B(n83), .Z(n280) );
  XOR2_X1 U247 ( .A(n278), .B(n280), .Z(product[14]) );
  NAND2_X1 U248 ( .A1(n14), .A2(n141), .ZN(n281) );
  NAND2_X1 U249 ( .A1(n141), .A2(n83), .ZN(n283) );
  BUF_X1 U250 ( .A(n234), .Z(n328) );
  XOR2_X1 U251 ( .A(n161), .B(n168), .Z(n284) );
  XOR2_X1 U252 ( .A(n120), .B(n284), .Z(n118) );
  NAND2_X1 U253 ( .A1(n120), .A2(n161), .ZN(n285) );
  NAND2_X1 U254 ( .A1(n120), .A2(n168), .ZN(n286) );
  NAND2_X1 U255 ( .A1(n161), .A2(n168), .ZN(n287) );
  NAND3_X1 U256 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n117) );
  NAND2_X1 U257 ( .A1(n332), .A2(n308), .ZN(n288) );
  CLKBUF_X1 U258 ( .A(n330), .Z(n289) );
  BUF_X2 U259 ( .A(n234), .Z(n330) );
  OR2_X1 U260 ( .A1(n114), .A2(n117), .ZN(n290) );
  BUF_X2 U261 ( .A(n225), .Z(n339) );
  XOR2_X1 U262 ( .A(n327), .B(a[2]), .Z(n291) );
  NAND2_X1 U263 ( .A1(n291), .A2(n227), .ZN(n292) );
  NAND2_X1 U264 ( .A1(n291), .A2(n227), .ZN(n293) );
  NAND2_X1 U265 ( .A1(n320), .A2(n227), .ZN(n223) );
  CLKBUF_X3 U266 ( .A(n236), .Z(n294) );
  BUF_X2 U267 ( .A(n216), .Z(n340) );
  BUF_X2 U268 ( .A(n235), .Z(n327) );
  CLKBUF_X1 U269 ( .A(n221), .Z(n295) );
  NAND2_X1 U270 ( .A1(n217), .A2(n225), .ZN(n221) );
  NAND2_X1 U271 ( .A1(n233), .A2(n297), .ZN(n298) );
  NAND2_X1 U272 ( .A1(n296), .A2(a[6]), .ZN(n299) );
  NAND2_X1 U273 ( .A1(n298), .A2(n299), .ZN(n217) );
  INV_X1 U274 ( .A(n233), .ZN(n296) );
  INV_X1 U275 ( .A(a[6]), .ZN(n297) );
  NAND2_X2 U276 ( .A1(n220), .A2(n244), .ZN(n224) );
  CLKBUF_X1 U277 ( .A(n276), .Z(n300) );
  CLKBUF_X1 U278 ( .A(n36), .Z(n301) );
  XNOR2_X1 U279 ( .A(n94), .B(n302), .ZN(n92) );
  XNOR2_X1 U280 ( .A(n97), .B(n144), .ZN(n302) );
  XNOR2_X1 U281 ( .A(n104), .B(n303), .ZN(n102) );
  XNOR2_X1 U282 ( .A(n109), .B(n106), .ZN(n303) );
  NAND2_X1 U283 ( .A1(n94), .A2(n97), .ZN(n304) );
  NAND2_X1 U284 ( .A1(n94), .A2(n144), .ZN(n305) );
  NAND2_X1 U285 ( .A1(n97), .A2(n144), .ZN(n306) );
  NAND3_X1 U286 ( .A1(n304), .A2(n305), .A3(n306), .ZN(n91) );
  OR2_X1 U287 ( .A1(n88), .A2(n91), .ZN(n323) );
  NAND2_X1 U288 ( .A1(n319), .A2(n226), .ZN(n307) );
  XOR2_X1 U289 ( .A(n330), .B(a[4]), .Z(n308) );
  NAND2_X1 U290 ( .A1(n308), .A2(n226), .ZN(n222) );
  AOI21_X1 U291 ( .B1(n322), .B2(n55), .A(n52), .ZN(n309) );
  AOI21_X1 U292 ( .B1(n322), .B2(n55), .A(n52), .ZN(n50) );
  CLKBUF_X1 U293 ( .A(n47), .Z(n310) );
  CLKBUF_X1 U294 ( .A(n29), .Z(n311) );
  OAI22_X1 U295 ( .A1(n293), .A2(n192), .B1(n191), .B2(n331), .ZN(n312) );
  CLKBUF_X1 U296 ( .A(n20), .Z(n313) );
  AOI21_X1 U297 ( .B1(n310), .B2(n39), .A(n40), .ZN(n314) );
  NAND2_X1 U298 ( .A1(n104), .A2(n109), .ZN(n315) );
  NAND2_X1 U299 ( .A1(n104), .A2(n106), .ZN(n316) );
  NAND2_X1 U300 ( .A1(n109), .A2(n106), .ZN(n317) );
  NAND3_X1 U301 ( .A1(n315), .A2(n316), .A3(n317), .ZN(n101) );
  NOR2_X1 U302 ( .A1(n102), .A2(n107), .ZN(n318) );
  OR2_X1 U303 ( .A1(n87), .A2(n86), .ZN(n324) );
  XOR2_X1 U304 ( .A(n330), .B(a[4]), .Z(n319) );
  XOR2_X1 U305 ( .A(n327), .B(a[2]), .Z(n320) );
  XNOR2_X1 U306 ( .A(n37), .B(n4), .ZN(product[9]) );
  INV_X1 U307 ( .A(n35), .ZN(n74) );
  INV_X1 U308 ( .A(n66), .ZN(n64) );
  INV_X1 U309 ( .A(n26), .ZN(n24) );
  NOR2_X1 U310 ( .A1(n102), .A2(n107), .ZN(n41) );
  INV_X1 U311 ( .A(n19), .ZN(n17) );
  NAND2_X1 U312 ( .A1(n324), .A2(n19), .ZN(n1) );
  XOR2_X1 U313 ( .A(n10), .B(n62), .Z(product[3]) );
  NAND2_X1 U314 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U315 ( .A(n60), .ZN(n80) );
  XOR2_X1 U316 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U317 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U318 ( .A(n56), .ZN(n79) );
  XOR2_X1 U319 ( .A(n32), .B(n3), .Z(product[10]) );
  AOI21_X1 U320 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U321 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U322 ( .A1(n76), .A2(n45), .ZN(n6) );
  INV_X1 U323 ( .A(n44), .ZN(n76) );
  XOR2_X1 U324 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U325 ( .A1(n323), .A2(n26), .ZN(n2) );
  XNOR2_X1 U326 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U327 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U328 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U329 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U330 ( .A1(n321), .A2(n66), .ZN(n11) );
  NAND2_X1 U331 ( .A1(n290), .A2(n49), .ZN(n7) );
  OR2_X1 U332 ( .A1(n171), .A2(n164), .ZN(n321) );
  XNOR2_X1 U333 ( .A(n158), .B(n146), .ZN(n106) );
  OR2_X1 U334 ( .A1(n158), .A2(n146), .ZN(n105) );
  NAND2_X1 U335 ( .A1(n108), .A2(n113), .ZN(n45) );
  NOR2_X1 U336 ( .A1(n122), .A2(n123), .ZN(n56) );
  NOR2_X1 U337 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U338 ( .A(n83), .ZN(n84) );
  OR2_X1 U339 ( .A1(n118), .A2(n121), .ZN(n322) );
  NAND2_X1 U340 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U341 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U342 ( .A1(n114), .A2(n117), .ZN(n49) );
  INV_X1 U343 ( .A(n69), .ZN(n67) );
  NAND2_X1 U344 ( .A1(n122), .A2(n123), .ZN(n57) );
  AND2_X1 U345 ( .A1(n340), .A2(n132), .ZN(n164) );
  OR2_X1 U346 ( .A1(n340), .A2(n231), .ZN(n199) );
  INV_X1 U347 ( .A(n128), .ZN(n149) );
  INV_X1 U348 ( .A(n89), .ZN(n90) );
  AND2_X1 U349 ( .A1(n340), .A2(n126), .ZN(n148) );
  OAI22_X1 U350 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  AND2_X1 U351 ( .A1(n340), .A2(n129), .ZN(n156) );
  OAI22_X1 U352 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U353 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI22_X1 U354 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OR2_X1 U355 ( .A1(n340), .A2(n230), .ZN(n190) );
  OAI22_X1 U356 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  BUF_X2 U357 ( .A(n227), .Z(n331) );
  BUF_X2 U358 ( .A(n226), .Z(n332) );
  INV_X1 U359 ( .A(n131), .ZN(n157) );
  INV_X1 U360 ( .A(n125), .ZN(n141) );
  OR2_X1 U361 ( .A1(n340), .A2(n229), .ZN(n181) );
  AND2_X1 U362 ( .A1(n274), .A2(n69), .ZN(product[1]) );
  OAI22_X1 U363 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U364 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  OR2_X1 U365 ( .A1(n340), .A2(n232), .ZN(n208) );
  AND2_X1 U366 ( .A1(n340), .A2(n135), .ZN(product[0]) );
  CLKBUF_X1 U367 ( .A(n234), .Z(n329) );
  XNOR2_X1 U368 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U369 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U370 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U371 ( .A(n233), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U372 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U373 ( .A(n340), .B(n233), .ZN(n180) );
  XNOR2_X1 U374 ( .A(n233), .B(b[1]), .ZN(n179) );
  INV_X1 U375 ( .A(n233), .ZN(n229) );
  XNOR2_X1 U376 ( .A(n236), .B(a[2]), .ZN(n227) );
  XNOR2_X1 U377 ( .A(n235), .B(a[4]), .ZN(n226) );
  NAND2_X1 U378 ( .A1(n73), .A2(n31), .ZN(n3) );
  NOR2_X1 U379 ( .A1(n92), .A2(n95), .ZN(n333) );
  NOR2_X1 U380 ( .A1(n92), .A2(n95), .ZN(n30) );
  XOR2_X1 U381 ( .A(n85), .B(n84), .Z(n334) );
  XOR2_X1 U382 ( .A(n300), .B(n334), .Z(product[13]) );
  NAND2_X1 U383 ( .A1(n276), .A2(n85), .ZN(n335) );
  NAND2_X1 U384 ( .A1(n276), .A2(n84), .ZN(n336) );
  NAND2_X1 U385 ( .A1(n85), .A2(n84), .ZN(n337) );
  NAND3_X1 U386 ( .A1(n335), .A2(n336), .A3(n337), .ZN(n14) );
  BUF_X2 U387 ( .A(n225), .Z(n338) );
  XNOR2_X1 U388 ( .A(n328), .B(a[6]), .ZN(n225) );
  NAND2_X1 U389 ( .A1(n74), .A2(n301), .ZN(n4) );
  INV_X1 U390 ( .A(n301), .ZN(n34) );
  NOR2_X1 U391 ( .A1(n96), .A2(n101), .ZN(n35) );
  INV_X1 U392 ( .A(n99), .ZN(n100) );
  INV_X1 U393 ( .A(n54), .ZN(n52) );
  NAND2_X1 U394 ( .A1(n322), .A2(n54), .ZN(n8) );
  INV_X1 U395 ( .A(n134), .ZN(n165) );
  NAND2_X1 U396 ( .A1(n124), .A2(n139), .ZN(n61) );
  NOR2_X1 U397 ( .A1(n124), .A2(n139), .ZN(n60) );
  NAND2_X1 U398 ( .A1(n96), .A2(n101), .ZN(n36) );
  NAND2_X1 U399 ( .A1(n92), .A2(n95), .ZN(n31) );
  OAI22_X1 U400 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  NAND2_X1 U401 ( .A1(n118), .A2(n121), .ZN(n54) );
  NAND2_X1 U402 ( .A1(n102), .A2(n107), .ZN(n42) );
  NAND2_X1 U403 ( .A1(n171), .A2(n164), .ZN(n66) );
  AOI21_X1 U404 ( .B1(n321), .B2(n67), .A(n64), .ZN(n62) );
  OAI21_X1 U405 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  INV_X1 U406 ( .A(n59), .ZN(n58) );
  OAI21_X1 U407 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  OAI22_X1 U408 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  XNOR2_X1 U409 ( .A(n233), .B(b[7]), .ZN(n173) );
  NAND2_X1 U410 ( .A1(n28), .A2(n323), .ZN(n21) );
  OAI21_X1 U411 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U412 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  XNOR2_X1 U413 ( .A(n327), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U414 ( .A(n326), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U415 ( .A(n327), .B(b[4]), .ZN(n194) );
  INV_X1 U416 ( .A(n326), .ZN(n231) );
  XNOR2_X1 U417 ( .A(n326), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U418 ( .A(n326), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U419 ( .A(n326), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U420 ( .A(n340), .B(n326), .ZN(n198) );
  XNOR2_X1 U421 ( .A(n327), .B(b[1]), .ZN(n197) );
  AOI21_X1 U422 ( .B1(n37), .B2(n277), .A(n311), .ZN(n27) );
  AOI21_X1 U423 ( .B1(n29), .B2(n323), .A(n24), .ZN(n22) );
  OAI21_X1 U424 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  NOR2_X1 U425 ( .A1(n35), .A2(n333), .ZN(n28) );
  INV_X1 U426 ( .A(n333), .ZN(n73) );
  XNOR2_X1 U427 ( .A(n8), .B(n55), .ZN(product[5]) );
  INV_X1 U428 ( .A(n310), .ZN(n46) );
  AOI21_X1 U429 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U430 ( .A1(n172), .A2(n140), .ZN(n69) );
  XNOR2_X1 U431 ( .A(n294), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U432 ( .A(n294), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U433 ( .A(n294), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U434 ( .A(n294), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U435 ( .A(n294), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U436 ( .A(n294), .B(b[3]), .ZN(n204) );
  XNOR2_X1 U437 ( .A(n340), .B(n294), .ZN(n207) );
  XNOR2_X1 U438 ( .A(n294), .B(b[1]), .ZN(n206) );
  INV_X1 U439 ( .A(n294), .ZN(n232) );
  XOR2_X1 U440 ( .A(n236), .B(n135), .Z(n220) );
  XOR2_X1 U441 ( .A(n7), .B(n309), .Z(product[6]) );
  OAI22_X1 U442 ( .A1(n182), .A2(n307), .B1(n182), .B2(n332), .ZN(n128) );
  OAI22_X1 U443 ( .A1(n307), .A2(n188), .B1(n187), .B2(n332), .ZN(n154) );
  OAI22_X1 U444 ( .A1(n307), .A2(n183), .B1(n182), .B2(n332), .ZN(n89) );
  OAI22_X1 U445 ( .A1(n307), .A2(n186), .B1(n185), .B2(n332), .ZN(n152) );
  OAI22_X1 U446 ( .A1(n222), .A2(n187), .B1(n186), .B2(n332), .ZN(n153) );
  OAI22_X1 U447 ( .A1(n307), .A2(n185), .B1(n184), .B2(n332), .ZN(n151) );
  OAI22_X1 U448 ( .A1(n307), .A2(n184), .B1(n183), .B2(n332), .ZN(n150) );
  INV_X1 U449 ( .A(n332), .ZN(n129) );
  OAI22_X1 U450 ( .A1(n288), .A2(n230), .B1(n190), .B2(n332), .ZN(n138) );
  OAI22_X1 U451 ( .A1(n288), .A2(n189), .B1(n188), .B2(n332), .ZN(n155) );
  INV_X1 U452 ( .A(n318), .ZN(n75) );
  OAI22_X1 U453 ( .A1(n173), .A2(n295), .B1(n173), .B2(n338), .ZN(n125) );
  OAI22_X1 U454 ( .A1(n295), .A2(n174), .B1(n173), .B2(n339), .ZN(n83) );
  NOR2_X1 U455 ( .A1(n318), .A2(n44), .ZN(n39) );
  OAI21_X1 U456 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI22_X1 U457 ( .A1(n295), .A2(n175), .B1(n174), .B2(n338), .ZN(n142) );
  OAI22_X1 U458 ( .A1(n295), .A2(n176), .B1(n175), .B2(n338), .ZN(n143) );
  OAI22_X1 U459 ( .A1(n295), .A2(n177), .B1(n176), .B2(n339), .ZN(n144) );
  XNOR2_X1 U460 ( .A(n329), .B(b[7]), .ZN(n182) );
  OAI22_X1 U461 ( .A1(n221), .A2(n178), .B1(n177), .B2(n339), .ZN(n145) );
  INV_X1 U462 ( .A(n339), .ZN(n126) );
  OAI22_X1 U463 ( .A1(n221), .A2(n179), .B1(n178), .B2(n338), .ZN(n146) );
  XNOR2_X1 U464 ( .A(n329), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U465 ( .A(n289), .B(b[5]), .ZN(n184) );
  OAI22_X1 U466 ( .A1(n221), .A2(n229), .B1(n181), .B2(n338), .ZN(n137) );
  OAI22_X1 U467 ( .A1(n221), .A2(n180), .B1(n179), .B2(n339), .ZN(n147) );
  XNOR2_X1 U468 ( .A(n289), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U469 ( .A(n329), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U470 ( .A(n329), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U471 ( .A(n340), .B(n330), .ZN(n189) );
  INV_X1 U472 ( .A(n329), .ZN(n230) );
  XNOR2_X1 U473 ( .A(n330), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U474 ( .A(n313), .B(n1), .ZN(product[12]) );
  INV_X1 U475 ( .A(n314), .ZN(n37) );
  AOI21_X1 U476 ( .B1(n20), .B2(n324), .A(n17), .ZN(n15) );
  OAI22_X1 U477 ( .A1(n292), .A2(n193), .B1(n192), .B2(n331), .ZN(n158) );
  OAI22_X1 U478 ( .A1(n293), .A2(n195), .B1(n194), .B2(n331), .ZN(n160) );
  OAI22_X1 U479 ( .A1(n223), .A2(n194), .B1(n193), .B2(n331), .ZN(n159) );
  OAI22_X1 U480 ( .A1(n293), .A2(n196), .B1(n195), .B2(n331), .ZN(n161) );
  OAI22_X1 U481 ( .A1(n292), .A2(n231), .B1(n199), .B2(n331), .ZN(n139) );
  OAI22_X1 U482 ( .A1(n292), .A2(n197), .B1(n196), .B2(n331), .ZN(n162) );
  OAI22_X1 U483 ( .A1(n223), .A2(n192), .B1(n191), .B2(n331), .ZN(n99) );
  OAI22_X1 U484 ( .A1(n191), .A2(n293), .B1(n191), .B2(n331), .ZN(n131) );
  INV_X1 U485 ( .A(n331), .ZN(n132) );
  OAI22_X1 U486 ( .A1(n223), .A2(n198), .B1(n197), .B2(n331), .ZN(n163) );
  INV_X2 U487 ( .A(n135), .ZN(n244) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n56,
         n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  FA_X1 U6 ( .A(A[11]), .B(B[11]), .CI(n17), .CO(n16), .S(SUM[11]) );
  AND2_X1 U86 ( .A1(A[1]), .A2(B[1]), .ZN(n129) );
  INV_X1 U87 ( .A(n129), .ZN(n56) );
  OR2_X1 U88 ( .A1(A[0]), .A2(B[0]), .ZN(n125) );
  CLKBUF_X1 U89 ( .A(n36), .Z(n126) );
  OR2_X2 U90 ( .A1(A[1]), .A2(B[1]), .ZN(n139) );
  AOI21_X1 U91 ( .B1(n41), .B2(n137), .A(n38), .ZN(n36) );
  AOI21_X1 U92 ( .B1(n139), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U93 ( .B1(n139), .B2(n128), .A(n129), .ZN(n52) );
  AND2_X1 U94 ( .A1(A[0]), .A2(B[0]), .ZN(n128) );
  CLKBUF_X1 U95 ( .A(n49), .Z(n130) );
  CLKBUF_X1 U96 ( .A(n33), .Z(n131) );
  CLKBUF_X1 U97 ( .A(n25), .Z(n132) );
  AOI21_X1 U98 ( .B1(n130), .B2(n138), .A(n46), .ZN(n133) );
  AOI21_X1 U99 ( .B1(n132), .B2(n140), .A(n22), .ZN(n134) );
  AOI21_X1 U100 ( .B1(n131), .B2(n141), .A(n30), .ZN(n135) );
  INV_X1 U101 ( .A(n24), .ZN(n22) );
  INV_X1 U102 ( .A(n40), .ZN(n38) );
  OAI21_X1 U103 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  AOI21_X1 U104 ( .B1(n49), .B2(n138), .A(n46), .ZN(n44) );
  INV_X1 U105 ( .A(n48), .ZN(n46) );
  AOI21_X1 U106 ( .B1(n33), .B2(n141), .A(n30), .ZN(n28) );
  INV_X1 U107 ( .A(n32), .ZN(n30) );
  NAND2_X1 U108 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U109 ( .A(n42), .ZN(n66) );
  NAND2_X1 U110 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U111 ( .A(n26), .ZN(n62) );
  NAND2_X1 U112 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U113 ( .A(n18), .ZN(n60) );
  NAND2_X1 U114 ( .A1(n138), .A2(n48), .ZN(n9) );
  NAND2_X1 U115 ( .A1(n141), .A2(n32), .ZN(n5) );
  NAND2_X1 U116 ( .A1(n140), .A2(n24), .ZN(n3) );
  XOR2_X1 U117 ( .A(n127), .B(n10), .Z(SUM[2]) );
  NAND2_X1 U118 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U119 ( .A(n50), .ZN(n68) );
  XOR2_X1 U120 ( .A(n126), .B(n6), .Z(SUM[6]) );
  NAND2_X1 U121 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U122 ( .A(n34), .ZN(n64) );
  XNOR2_X1 U123 ( .A(n41), .B(n7), .ZN(SUM[5]) );
  NAND2_X1 U124 ( .A1(n137), .A2(n40), .ZN(n7) );
  XNOR2_X1 U125 ( .A(n11), .B(n128), .ZN(SUM[1]) );
  NAND2_X1 U126 ( .A1(n139), .A2(n56), .ZN(n11) );
  XNOR2_X1 U127 ( .A(n13), .B(n136), .ZN(SUM[15]) );
  XNOR2_X1 U128 ( .A(B[15]), .B(A[15]), .ZN(n136) );
  NOR2_X1 U129 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  OR2_X1 U130 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  OR2_X1 U131 ( .A1(A[3]), .A2(B[3]), .ZN(n138) );
  NOR2_X1 U132 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U133 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U134 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U135 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U136 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U137 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U138 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U139 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  NAND2_X1 U140 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  OR2_X1 U141 ( .A1(A[9]), .A2(B[9]), .ZN(n140) );
  OR2_X1 U142 ( .A1(A[7]), .A2(B[7]), .ZN(n141) );
  NAND2_X1 U143 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U144 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U145 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U146 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  AND2_X1 U147 ( .A1(n125), .A2(n59), .ZN(SUM[0]) );
  OAI21_X1 U148 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U149 ( .A(n131), .B(n5), .ZN(SUM[7]) );
  XNOR2_X1 U150 ( .A(n132), .B(n3), .ZN(SUM[9]) );
  XOR2_X1 U151 ( .A(n133), .B(n8), .Z(SUM[4]) );
  AOI21_X1 U152 ( .B1(n25), .B2(n140), .A(n22), .ZN(n20) );
  NAND2_X1 U153 ( .A1(A[0]), .A2(B[0]), .ZN(n59) );
  XOR2_X1 U154 ( .A(n134), .B(n2), .Z(SUM[10]) );
  XNOR2_X1 U155 ( .A(n130), .B(n9), .ZN(SUM[3]) );
  XOR2_X1 U156 ( .A(n135), .B(n4), .Z(SUM[8]) );
  OAI21_X1 U157 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U158 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X1 U159 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
endmodule


module add_layer_WIDTH16_0 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_0_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_11_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n56,
         n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n137, n138, n139, n140, n141, n142,
         n143;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  FA_X1 U6 ( .A(A[11]), .B(B[11]), .CI(n17), .CO(n16), .S(SUM[11]) );
  CLKBUF_X1 U86 ( .A(n36), .Z(n125) );
  AOI21_X1 U87 ( .B1(n41), .B2(n141), .A(n38), .ZN(n36) );
  OR2_X1 U88 ( .A1(A[0]), .A2(B[0]), .ZN(n126) );
  AND2_X1 U89 ( .A1(A[1]), .A2(B[1]), .ZN(n129) );
  INV_X1 U90 ( .A(n129), .ZN(n56) );
  OR2_X2 U91 ( .A1(A[1]), .A2(B[1]), .ZN(n140) );
  AOI21_X1 U92 ( .B1(n140), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U93 ( .B1(n140), .B2(n128), .A(n129), .ZN(n52) );
  AND2_X1 U94 ( .A1(A[0]), .A2(B[0]), .ZN(n128) );
  CLKBUF_X1 U95 ( .A(n25), .Z(n130) );
  CLKBUF_X1 U96 ( .A(n41), .Z(n131) );
  AOI21_X1 U97 ( .B1(n130), .B2(n142), .A(n22), .ZN(n132) );
  CLKBUF_X1 U98 ( .A(n33), .Z(n133) );
  AOI21_X1 U99 ( .B1(n135), .B2(n139), .A(n46), .ZN(n134) );
  CLKBUF_X1 U100 ( .A(n49), .Z(n135) );
  AOI21_X1 U101 ( .B1(n49), .B2(n139), .A(n46), .ZN(n44) );
  AND2_X1 U102 ( .A1(n126), .A2(n59), .ZN(SUM[0]) );
  INV_X1 U103 ( .A(n40), .ZN(n38) );
  AOI21_X1 U104 ( .B1(n25), .B2(n142), .A(n22), .ZN(n20) );
  INV_X1 U105 ( .A(n24), .ZN(n22) );
  INV_X1 U106 ( .A(n48), .ZN(n46) );
  NAND2_X1 U107 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U108 ( .A(n34), .ZN(n64) );
  NAND2_X1 U109 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U110 ( .A(n26), .ZN(n62) );
  NAND2_X1 U111 ( .A1(n138), .A2(n32), .ZN(n5) );
  XOR2_X1 U112 ( .A(n132), .B(n2), .Z(SUM[10]) );
  NAND2_X1 U113 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U114 ( .A(n18), .ZN(n60) );
  XOR2_X1 U115 ( .A(n127), .B(n10), .Z(SUM[2]) );
  NAND2_X1 U116 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U117 ( .A(n50), .ZN(n68) );
  XOR2_X1 U118 ( .A(n134), .B(n8), .Z(SUM[4]) );
  NAND2_X1 U119 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U120 ( .A(n42), .ZN(n66) );
  XNOR2_X1 U121 ( .A(n135), .B(n9), .ZN(SUM[3]) );
  NAND2_X1 U122 ( .A1(n139), .A2(n48), .ZN(n9) );
  XNOR2_X1 U123 ( .A(n130), .B(n3), .ZN(SUM[9]) );
  NAND2_X1 U124 ( .A1(n142), .A2(n24), .ZN(n3) );
  XNOR2_X1 U125 ( .A(n131), .B(n7), .ZN(SUM[5]) );
  NAND2_X1 U126 ( .A1(n141), .A2(n40), .ZN(n7) );
  XNOR2_X1 U127 ( .A(n11), .B(n128), .ZN(SUM[1]) );
  NAND2_X1 U128 ( .A1(n140), .A2(n56), .ZN(n11) );
  INV_X1 U129 ( .A(n32), .ZN(n30) );
  XNOR2_X1 U130 ( .A(n13), .B(n137), .ZN(SUM[15]) );
  XNOR2_X1 U131 ( .A(B[15]), .B(A[15]), .ZN(n137) );
  OR2_X1 U132 ( .A1(A[7]), .A2(B[7]), .ZN(n138) );
  OR2_X1 U133 ( .A1(A[3]), .A2(B[3]), .ZN(n139) );
  NOR2_X1 U134 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  NOR2_X1 U135 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U136 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U137 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U138 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U140 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U141 ( .A1(A[0]), .A2(B[0]), .ZN(n59) );
  NAND2_X1 U142 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U143 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  OR2_X1 U144 ( .A1(A[5]), .A2(B[5]), .ZN(n141) );
  OR2_X1 U145 ( .A1(A[9]), .A2(B[9]), .ZN(n142) );
  NAND2_X1 U146 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  NAND2_X1 U147 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U148 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U149 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U150 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  OAI21_X1 U151 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  OAI21_X1 U152 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  AOI21_X1 U153 ( .B1(n133), .B2(n138), .A(n30), .ZN(n143) );
  AOI21_X1 U154 ( .B1(n33), .B2(n138), .A(n30), .ZN(n28) );
  XNOR2_X1 U155 ( .A(n133), .B(n5), .ZN(SUM[7]) );
  OAI21_X1 U156 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  XOR2_X1 U157 ( .A(n125), .B(n6), .Z(SUM[6]) );
  OAI21_X1 U158 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U159 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U160 ( .A(n143), .B(n4), .Z(SUM[8]) );
endmodule


module add_layer_WIDTH16_11 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_11_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n21,
         n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37, n38, n39,
         n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55, n56, n57,
         n61, n62, n64, n65, n67, n69, n71, n73, n75, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173;

  NAND2_X1 U94 ( .A1(A[13]), .A2(B[13]), .ZN(n149) );
  AOI21_X1 U95 ( .B1(n46), .B2(n168), .A(n43), .ZN(n41) );
  AND2_X1 U96 ( .A1(n170), .A2(n64), .ZN(SUM[0]) );
  NAND3_X1 U97 ( .A1(n138), .A2(n137), .A3(n139), .ZN(n133) );
  OAI21_X1 U98 ( .B1(n142), .B2(n141), .A(n21), .ZN(n134) );
  OAI21_X1 U99 ( .B1(n142), .B2(n141), .A(n21), .ZN(n135) );
  OAI21_X1 U100 ( .B1(n142), .B2(n141), .A(n21), .ZN(n65) );
  XOR2_X1 U101 ( .A(A[12]), .B(B[12]), .Z(n136) );
  XOR2_X1 U102 ( .A(n135), .B(n136), .Z(SUM[12]) );
  NAND2_X1 U103 ( .A1(n65), .A2(A[12]), .ZN(n137) );
  NAND2_X1 U104 ( .A1(n134), .A2(B[12]), .ZN(n138) );
  NAND2_X1 U105 ( .A1(A[12]), .A2(B[12]), .ZN(n139) );
  NAND3_X1 U106 ( .A1(n138), .A2(n137), .A3(n139), .ZN(n16) );
  CLKBUF_X1 U107 ( .A(n133), .Z(n140) );
  INV_X1 U108 ( .A(n172), .ZN(n141) );
  INV_X1 U109 ( .A(n22), .ZN(n142) );
  AOI21_X1 U110 ( .B1(n54), .B2(n167), .A(n51), .ZN(n143) );
  AOI21_X1 U111 ( .B1(n54), .B2(n167), .A(n51), .ZN(n49) );
  CLKBUF_X1 U112 ( .A(n46), .Z(n144) );
  CLKBUF_X1 U113 ( .A(n54), .Z(n145) );
  NAND3_X1 U114 ( .A1(n151), .A2(n150), .A3(n149), .ZN(n146) );
  NAND3_X1 U115 ( .A1(n151), .A2(n150), .A3(n149), .ZN(n147) );
  XOR2_X1 U116 ( .A(A[13]), .B(B[13]), .Z(n148) );
  XOR2_X1 U117 ( .A(n148), .B(n140), .Z(SUM[13]) );
  NAND2_X1 U118 ( .A1(A[13]), .A2(n16), .ZN(n150) );
  NAND2_X1 U119 ( .A1(B[13]), .A2(n133), .ZN(n151) );
  NAND3_X1 U120 ( .A1(n151), .A2(n150), .A3(n149), .ZN(n15) );
  XOR2_X1 U121 ( .A(A[14]), .B(B[14]), .Z(n152) );
  XOR2_X1 U122 ( .A(n152), .B(n147), .Z(SUM[14]) );
  NAND2_X1 U123 ( .A1(A[14]), .A2(B[14]), .ZN(n153) );
  NAND2_X1 U124 ( .A1(n15), .A2(A[14]), .ZN(n154) );
  NAND2_X1 U125 ( .A1(B[14]), .A2(n146), .ZN(n155) );
  NAND3_X1 U126 ( .A1(n155), .A2(n154), .A3(n153), .ZN(n14) );
  OR2_X1 U127 ( .A1(A[1]), .A2(B[1]), .ZN(n156) );
  INV_X1 U128 ( .A(n61), .ZN(n157) );
  OR2_X1 U129 ( .A1(A[1]), .A2(B[1]), .ZN(n169) );
  AND2_X1 U130 ( .A1(A[1]), .A2(B[1]), .ZN(n160) );
  INV_X1 U131 ( .A(n160), .ZN(n61) );
  AND2_X1 U132 ( .A1(A[0]), .A2(B[0]), .ZN(n158) );
  CLKBUF_X1 U133 ( .A(n30), .Z(n159) );
  AOI21_X1 U134 ( .B1(n159), .B2(n171), .A(n27), .ZN(n161) );
  CLKBUF_X1 U135 ( .A(n38), .Z(n162) );
  CLKBUF_X1 U136 ( .A(n22), .Z(n163) );
  AOI21_X1 U137 ( .B1(n38), .B2(n173), .A(n35), .ZN(n164) );
  AOI21_X1 U138 ( .B1(n169), .B2(n158), .A(n160), .ZN(n165) );
  INV_X1 U139 ( .A(n29), .ZN(n27) );
  AOI21_X1 U140 ( .B1(n156), .B2(n62), .A(n157), .ZN(n57) );
  OAI21_X1 U141 ( .B1(n165), .B2(n55), .A(n56), .ZN(n54) );
  INV_X1 U142 ( .A(n53), .ZN(n51) );
  INV_X1 U143 ( .A(n45), .ZN(n43) );
  AOI21_X1 U144 ( .B1(n162), .B2(n173), .A(n35), .ZN(n33) );
  INV_X1 U145 ( .A(n37), .ZN(n35) );
  NAND2_X1 U146 ( .A1(n67), .A2(n24), .ZN(n3) );
  INV_X1 U147 ( .A(n23), .ZN(n67) );
  NAND2_X1 U148 ( .A1(n71), .A2(n40), .ZN(n7) );
  INV_X1 U149 ( .A(n39), .ZN(n71) );
  NAND2_X1 U150 ( .A1(n69), .A2(n32), .ZN(n5) );
  INV_X1 U151 ( .A(n31), .ZN(n69) );
  NAND2_X1 U152 ( .A1(n172), .A2(n21), .ZN(n2) );
  NAND2_X1 U153 ( .A1(n168), .A2(n45), .ZN(n8) );
  NAND2_X1 U154 ( .A1(n173), .A2(n37), .ZN(n6) );
  NAND2_X1 U155 ( .A1(n171), .A2(n29), .ZN(n4) );
  NAND2_X1 U156 ( .A1(n167), .A2(n53), .ZN(n10) );
  XNOR2_X1 U157 ( .A(n12), .B(n62), .ZN(SUM[1]) );
  NAND2_X1 U158 ( .A1(n156), .A2(n61), .ZN(n12) );
  NAND2_X1 U159 ( .A1(n75), .A2(n56), .ZN(n11) );
  INV_X1 U160 ( .A(n55), .ZN(n75) );
  NAND2_X1 U161 ( .A1(n73), .A2(n48), .ZN(n9) );
  INV_X1 U162 ( .A(n47), .ZN(n73) );
  XNOR2_X1 U163 ( .A(n14), .B(n166), .ZN(SUM[15]) );
  XNOR2_X1 U164 ( .A(B[15]), .B(A[15]), .ZN(n166) );
  NOR2_X1 U165 ( .A1(A[2]), .A2(B[2]), .ZN(n55) );
  OR2_X1 U166 ( .A1(A[3]), .A2(B[3]), .ZN(n167) );
  OR2_X1 U167 ( .A1(A[5]), .A2(B[5]), .ZN(n168) );
  NOR2_X1 U168 ( .A1(A[6]), .A2(B[6]), .ZN(n39) );
  NOR2_X1 U169 ( .A1(A[8]), .A2(B[8]), .ZN(n31) );
  NOR2_X1 U170 ( .A1(A[4]), .A2(B[4]), .ZN(n47) );
  NOR2_X1 U171 ( .A1(A[10]), .A2(B[10]), .ZN(n23) );
  OR2_X1 U172 ( .A1(A[0]), .A2(B[0]), .ZN(n170) );
  NAND2_X1 U173 ( .A1(A[9]), .A2(B[9]), .ZN(n29) );
  NAND2_X1 U174 ( .A1(A[7]), .A2(B[7]), .ZN(n37) );
  NAND2_X1 U175 ( .A1(A[3]), .A2(B[3]), .ZN(n53) );
  NAND2_X1 U176 ( .A1(A[5]), .A2(B[5]), .ZN(n45) );
  NAND2_X1 U177 ( .A1(A[11]), .A2(B[11]), .ZN(n21) );
  NAND2_X1 U178 ( .A1(A[2]), .A2(B[2]), .ZN(n56) );
  OR2_X1 U179 ( .A1(A[9]), .A2(B[9]), .ZN(n171) );
  OR2_X1 U180 ( .A1(A[11]), .A2(B[11]), .ZN(n172) );
  OR2_X1 U181 ( .A1(A[7]), .A2(B[7]), .ZN(n173) );
  NAND2_X1 U182 ( .A1(A[6]), .A2(B[6]), .ZN(n40) );
  NAND2_X1 U183 ( .A1(A[8]), .A2(B[8]), .ZN(n32) );
  NAND2_X1 U184 ( .A1(A[4]), .A2(B[4]), .ZN(n48) );
  NAND2_X1 U185 ( .A1(A[10]), .A2(B[10]), .ZN(n24) );
  XNOR2_X1 U186 ( .A(n159), .B(n4), .ZN(SUM[9]) );
  XNOR2_X1 U187 ( .A(n144), .B(n8), .ZN(SUM[5]) );
  XOR2_X1 U188 ( .A(n143), .B(n9), .Z(SUM[4]) );
  OAI21_X1 U189 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  INV_X1 U190 ( .A(n64), .ZN(n62) );
  XNOR2_X1 U191 ( .A(n145), .B(n10), .ZN(SUM[3]) );
  XOR2_X1 U192 ( .A(n41), .B(n7), .Z(SUM[6]) );
  NAND2_X1 U193 ( .A1(A[0]), .A2(B[0]), .ZN(n64) );
  AOI21_X1 U194 ( .B1(n30), .B2(n171), .A(n27), .ZN(n25) );
  XNOR2_X1 U195 ( .A(n162), .B(n6), .ZN(SUM[7]) );
  OAI21_X1 U196 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  XOR2_X1 U197 ( .A(n57), .B(n11), .Z(SUM[2]) );
  XOR2_X1 U198 ( .A(n33), .B(n5), .Z(SUM[8]) );
  OAI21_X1 U199 ( .B1(n164), .B2(n31), .A(n32), .ZN(n30) );
  XNOR2_X1 U200 ( .A(n163), .B(n2), .ZN(SUM[11]) );
  OAI21_X1 U201 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
  XOR2_X1 U202 ( .A(n161), .B(n3), .Z(SUM[10]) );
endmodule


module add_layer_WIDTH16_4 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_4_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_0 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_4 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_0 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_0 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_11 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_0 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_0 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0 \genblk1[0].mult  ( .clk(clk), .ia(
        {\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15 \genblk1[1].mult  ( .clk(clk), 
        .ia({\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14 \genblk1[2].mult  ( .clk(clk), 
        .ia({\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13 \genblk1[3].mult  ( .clk(clk), 
        .ia({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_0 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n31, n32, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n74,
         n75, n76, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n128,
         n131, n132, n134, n135, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n216,
         n217, n219, n220, n221, n222, n223, n224, n225, n227, n229, n230,
         n231, n232, n233, n234, n235, n236, n244, n274, n275, n276, n277,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n342, n343, n344, n345,
         n346, n347, n348;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n150), .B(n326), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n145), .B(n100), .CI(n151), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n159), .B(n153), .CI(n166), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n160), .B(n148), .CI(n167), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n138), .B(n155), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  OR2_X1 U237 ( .A1(n319), .A2(n95), .ZN(n274) );
  OR2_X1 U238 ( .A1(n172), .A2(n140), .ZN(n275) );
  CLKBUF_X1 U239 ( .A(n235), .Z(n276) );
  CLKBUF_X1 U240 ( .A(n235), .Z(n277) );
  CLKBUF_X1 U241 ( .A(n216), .Z(n348) );
  CLKBUF_X1 U242 ( .A(n216), .Z(n289) );
  AND3_X1 U243 ( .A1(n315), .A2(n314), .A3(n313), .ZN(product[15]) );
  XNOR2_X1 U244 ( .A(n279), .B(n296), .ZN(product[14]) );
  XNOR2_X1 U245 ( .A(n141), .B(n83), .ZN(n279) );
  OR2_X1 U246 ( .A1(n114), .A2(n117), .ZN(n280) );
  INV_X1 U247 ( .A(n74), .ZN(n281) );
  XNOR2_X1 U248 ( .A(n234), .B(a[4]), .ZN(n282) );
  INV_X1 U249 ( .A(n230), .ZN(n283) );
  XOR2_X1 U250 ( .A(n235), .B(a[4]), .Z(n284) );
  XOR2_X1 U251 ( .A(n233), .B(a[6]), .Z(n285) );
  XOR2_X1 U252 ( .A(n233), .B(a[6]), .Z(n286) );
  XNOR2_X1 U253 ( .A(n234), .B(a[6]), .ZN(n287) );
  XNOR2_X1 U254 ( .A(n234), .B(a[6]), .ZN(n288) );
  XNOR2_X1 U255 ( .A(n234), .B(a[6]), .ZN(n225) );
  CLKBUF_X1 U256 ( .A(n50), .Z(n290) );
  CLKBUF_X1 U257 ( .A(n236), .Z(n291) );
  NOR2_X1 U258 ( .A1(n281), .A2(n333), .ZN(n292) );
  NAND2_X1 U259 ( .A1(n219), .A2(n347), .ZN(n293) );
  CLKBUF_X1 U260 ( .A(n235), .Z(n294) );
  NAND3_X1 U261 ( .A1(n312), .A2(n311), .A3(n310), .ZN(n295) );
  NAND3_X1 U262 ( .A1(n311), .A2(n310), .A3(n312), .ZN(n296) );
  CLKBUF_X1 U263 ( .A(n70), .Z(n297) );
  CLKBUF_X1 U264 ( .A(n345), .Z(n298) );
  XNOR2_X2 U265 ( .A(n236), .B(a[2]), .ZN(n299) );
  CLKBUF_X1 U266 ( .A(n40), .Z(n300) );
  NAND2_X1 U267 ( .A1(n235), .A2(n302), .ZN(n303) );
  NAND2_X1 U268 ( .A1(n301), .A2(a[2]), .ZN(n304) );
  NAND2_X1 U269 ( .A1(n303), .A2(n304), .ZN(n219) );
  INV_X1 U270 ( .A(n235), .ZN(n301) );
  INV_X1 U271 ( .A(a[2]), .ZN(n302) );
  BUF_X1 U272 ( .A(n219), .Z(n325) );
  XNOR2_X2 U273 ( .A(n235), .B(a[4]), .ZN(n342) );
  AOI21_X1 U274 ( .B1(n340), .B2(n55), .A(n52), .ZN(n50) );
  NAND2_X1 U275 ( .A1(n236), .A2(n306), .ZN(n307) );
  NAND2_X1 U276 ( .A1(n305), .A2(n135), .ZN(n308) );
  NAND2_X1 U277 ( .A1(n307), .A2(n308), .ZN(n220) );
  INV_X1 U278 ( .A(n236), .ZN(n305) );
  INV_X1 U279 ( .A(n135), .ZN(n306) );
  XOR2_X1 U280 ( .A(n85), .B(n84), .Z(n309) );
  XOR2_X1 U281 ( .A(n309), .B(n297), .Z(product[13]) );
  NAND2_X1 U282 ( .A1(n85), .A2(n84), .ZN(n310) );
  NAND2_X1 U283 ( .A1(n70), .A2(n85), .ZN(n311) );
  NAND2_X1 U284 ( .A1(n84), .A2(n70), .ZN(n312) );
  NAND3_X1 U285 ( .A1(n312), .A2(n311), .A3(n310), .ZN(n14) );
  NAND2_X1 U286 ( .A1(n141), .A2(n83), .ZN(n313) );
  NAND2_X1 U287 ( .A1(n141), .A2(n14), .ZN(n314) );
  NAND2_X1 U288 ( .A1(n83), .A2(n295), .ZN(n315) );
  OR2_X2 U289 ( .A1(n282), .A2(n284), .ZN(n316) );
  NOR2_X2 U290 ( .A1(n108), .A2(n113), .ZN(n44) );
  XNOR2_X1 U291 ( .A(n104), .B(n317), .ZN(n102) );
  XNOR2_X1 U292 ( .A(n109), .B(n106), .ZN(n317) );
  CLKBUF_X1 U293 ( .A(n36), .Z(n318) );
  CLKBUF_X1 U294 ( .A(n92), .Z(n319) );
  OR2_X2 U295 ( .A1(n320), .A2(n321), .ZN(n222) );
  XNOR2_X1 U296 ( .A(n234), .B(a[4]), .ZN(n320) );
  XOR2_X1 U297 ( .A(n235), .B(a[4]), .Z(n321) );
  CLKBUF_X1 U298 ( .A(n20), .Z(n322) );
  CLKBUF_X1 U299 ( .A(n47), .Z(n323) );
  CLKBUF_X1 U300 ( .A(n29), .Z(n324) );
  OAI22_X1 U301 ( .A1(n345), .A2(n192), .B1(n191), .B2(n299), .ZN(n326) );
  NAND2_X1 U302 ( .A1(n104), .A2(n109), .ZN(n327) );
  NAND2_X1 U303 ( .A1(n104), .A2(n106), .ZN(n328) );
  NAND2_X1 U304 ( .A1(n109), .A2(n106), .ZN(n329) );
  NAND3_X1 U305 ( .A1(n327), .A2(n328), .A3(n329), .ZN(n101) );
  AOI21_X1 U306 ( .B1(n39), .B2(n323), .A(n300), .ZN(n330) );
  CLKBUF_X1 U307 ( .A(n287), .Z(n331) );
  NOR2_X1 U308 ( .A1(n92), .A2(n95), .ZN(n332) );
  NOR2_X1 U309 ( .A1(n92), .A2(n95), .ZN(n333) );
  NOR2_X1 U310 ( .A1(n102), .A2(n107), .ZN(n334) );
  NAND2_X1 U311 ( .A1(n220), .A2(n244), .ZN(n335) );
  NAND2_X1 U312 ( .A1(n220), .A2(n244), .ZN(n336) );
  INV_X1 U313 ( .A(n35), .ZN(n74) );
  INV_X1 U314 ( .A(n323), .ZN(n46) );
  XNOR2_X1 U315 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U316 ( .A1(n74), .A2(n318), .ZN(n4) );
  INV_X1 U317 ( .A(n318), .ZN(n34) );
  INV_X1 U318 ( .A(n26), .ZN(n24) );
  OAI21_X1 U319 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  NAND2_X1 U320 ( .A1(n280), .A2(n49), .ZN(n7) );
  NAND2_X1 U321 ( .A1(n339), .A2(n19), .ZN(n1) );
  XOR2_X1 U322 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U323 ( .A1(n76), .A2(n45), .ZN(n6) );
  INV_X1 U324 ( .A(n44), .ZN(n76) );
  XOR2_X1 U325 ( .A(n10), .B(n62), .Z(product[3]) );
  NAND2_X1 U326 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U327 ( .A(n60), .ZN(n80) );
  XOR2_X1 U328 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U329 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U330 ( .A(n56), .ZN(n79) );
  XOR2_X1 U331 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U332 ( .A1(n274), .A2(n31), .ZN(n3) );
  AOI21_X1 U333 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U334 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U335 ( .A1(n338), .A2(n26), .ZN(n2) );
  NOR2_X1 U336 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U337 ( .A1(n96), .A2(n101), .ZN(n36) );
  XNOR2_X1 U338 ( .A(n8), .B(n55), .ZN(product[5]) );
  XNOR2_X1 U339 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U340 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U341 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U342 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U343 ( .A1(n337), .A2(n66), .ZN(n11) );
  INV_X1 U344 ( .A(n19), .ZN(n17) );
  OR2_X1 U345 ( .A1(n158), .A2(n146), .ZN(n105) );
  NOR2_X1 U346 ( .A1(n102), .A2(n107), .ZN(n41) );
  XNOR2_X1 U347 ( .A(n158), .B(n146), .ZN(n106) );
  NOR2_X1 U348 ( .A1(n122), .A2(n123), .ZN(n56) );
  OR2_X1 U349 ( .A1(n171), .A2(n164), .ZN(n337) );
  NAND2_X1 U350 ( .A1(n108), .A2(n113), .ZN(n45) );
  NOR2_X1 U351 ( .A1(n114), .A2(n117), .ZN(n48) );
  NAND2_X1 U352 ( .A1(n102), .A2(n107), .ZN(n42) );
  NOR2_X1 U353 ( .A1(n124), .A2(n139), .ZN(n60) );
  INV_X1 U354 ( .A(n83), .ZN(n84) );
  OR2_X1 U355 ( .A1(n88), .A2(n91), .ZN(n338) );
  NAND2_X1 U356 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U357 ( .A1(n87), .A2(n86), .ZN(n19) );
  INV_X1 U358 ( .A(n69), .ZN(n67) );
  NAND2_X1 U359 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U360 ( .A1(n122), .A2(n123), .ZN(n57) );
  OR2_X1 U361 ( .A1(n87), .A2(n86), .ZN(n339) );
  NAND2_X1 U362 ( .A1(n92), .A2(n95), .ZN(n31) );
  OR2_X1 U363 ( .A1(n118), .A2(n121), .ZN(n340) );
  OR2_X1 U364 ( .A1(n289), .A2(n231), .ZN(n199) );
  INV_X1 U365 ( .A(n128), .ZN(n149) );
  INV_X1 U366 ( .A(n89), .ZN(n90) );
  AND2_X1 U367 ( .A1(n289), .A2(n284), .ZN(n156) );
  OAI22_X1 U368 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OR2_X1 U369 ( .A1(n348), .A2(n230), .ZN(n190) );
  AND2_X1 U370 ( .A1(n289), .A2(n126), .ZN(n148) );
  INV_X1 U371 ( .A(n125), .ZN(n141) );
  AND2_X1 U372 ( .A1(n275), .A2(n69), .ZN(product[1]) );
  AND2_X1 U373 ( .A1(n289), .A2(n132), .ZN(n164) );
  OR2_X1 U374 ( .A1(n348), .A2(n229), .ZN(n181) );
  INV_X1 U375 ( .A(n135), .ZN(n244) );
  OAI22_X1 U376 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  OR2_X1 U377 ( .A1(n289), .A2(n232), .ZN(n208) );
  NAND2_X1 U378 ( .A1(n220), .A2(n244), .ZN(n224) );
  AND2_X1 U379 ( .A1(n289), .A2(n135), .ZN(product[0]) );
  NAND2_X1 U380 ( .A1(n219), .A2(n227), .ZN(n345) );
  NAND2_X1 U381 ( .A1(n219), .A2(n347), .ZN(n346) );
  XNOR2_X1 U382 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U383 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U384 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U385 ( .A(n348), .B(n233), .ZN(n180) );
  INV_X1 U386 ( .A(n233), .ZN(n229) );
  INV_X1 U387 ( .A(n99), .ZN(n100) );
  NAND2_X1 U388 ( .A1(n171), .A2(n164), .ZN(n66) );
  NAND2_X1 U389 ( .A1(n124), .A2(n139), .ZN(n61) );
  OAI22_X1 U390 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U391 ( .A1(n336), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  XNOR2_X1 U392 ( .A(n233), .B(b[6]), .ZN(n174) );
  INV_X1 U393 ( .A(n131), .ZN(n157) );
  NAND2_X1 U394 ( .A1(n217), .A2(n225), .ZN(n343) );
  NAND2_X1 U395 ( .A1(n286), .A2(n287), .ZN(n344) );
  NAND2_X1 U396 ( .A1(n285), .A2(n288), .ZN(n221) );
  XOR2_X1 U397 ( .A(n233), .B(a[6]), .Z(n217) );
  INV_X1 U398 ( .A(n54), .ZN(n52) );
  NAND2_X1 U399 ( .A1(n340), .A2(n54), .ZN(n8) );
  XNOR2_X1 U400 ( .A(n233), .B(b[7]), .ZN(n173) );
  OAI22_X1 U401 ( .A1(n336), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  NAND2_X1 U402 ( .A1(n172), .A2(n140), .ZN(n69) );
  OAI21_X1 U403 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  INV_X1 U404 ( .A(n234), .ZN(n230) );
  XNOR2_X1 U405 ( .A(n283), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U406 ( .A(n234), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U407 ( .A(n234), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U408 ( .A(n283), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U409 ( .A(n234), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U410 ( .A(n348), .B(n234), .ZN(n189) );
  INV_X1 U411 ( .A(n134), .ZN(n165) );
  OAI22_X1 U412 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  OAI22_X1 U413 ( .A1(n335), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  XNOR2_X1 U414 ( .A(n236), .B(a[2]), .ZN(n347) );
  NAND2_X1 U415 ( .A1(n325), .A2(n227), .ZN(n223) );
  XNOR2_X1 U416 ( .A(n236), .B(a[2]), .ZN(n227) );
  NAND2_X1 U417 ( .A1(n28), .A2(n338), .ZN(n21) );
  NOR2_X1 U418 ( .A1(n35), .A2(n333), .ZN(n28) );
  AOI21_X1 U419 ( .B1(n29), .B2(n338), .A(n24), .ZN(n22) );
  AOI21_X1 U420 ( .B1(n37), .B2(n292), .A(n324), .ZN(n27) );
  OAI21_X1 U421 ( .B1(n332), .B2(n36), .A(n31), .ZN(n29) );
  INV_X1 U422 ( .A(n59), .ZN(n58) );
  AOI21_X1 U423 ( .B1(n337), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U424 ( .A(n66), .ZN(n64) );
  OAI22_X1 U425 ( .A1(n336), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  NAND2_X1 U426 ( .A1(n118), .A2(n121), .ZN(n54) );
  OAI22_X1 U427 ( .A1(n182), .A2(n316), .B1(n182), .B2(n342), .ZN(n128) );
  OAI22_X1 U428 ( .A1(n316), .A2(n188), .B1(n187), .B2(n342), .ZN(n154) );
  OAI22_X1 U429 ( .A1(n316), .A2(n183), .B1(n182), .B2(n342), .ZN(n89) );
  OAI22_X1 U430 ( .A1(n222), .A2(n187), .B1(n186), .B2(n342), .ZN(n153) );
  OAI22_X1 U431 ( .A1(n316), .A2(n186), .B1(n185), .B2(n342), .ZN(n152) );
  OAI22_X1 U432 ( .A1(n316), .A2(n185), .B1(n184), .B2(n342), .ZN(n151) );
  OAI22_X1 U433 ( .A1(n316), .A2(n184), .B1(n183), .B2(n342), .ZN(n150) );
  XNOR2_X1 U434 ( .A(n276), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U435 ( .A(n277), .B(b[4]), .ZN(n194) );
  OAI22_X1 U436 ( .A1(n222), .A2(n230), .B1(n190), .B2(n342), .ZN(n138) );
  OAI22_X1 U437 ( .A1(n222), .A2(n189), .B1(n188), .B2(n342), .ZN(n155) );
  INV_X1 U438 ( .A(n294), .ZN(n231) );
  XNOR2_X1 U439 ( .A(n294), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U440 ( .A(n289), .B(n294), .ZN(n198) );
  XNOR2_X1 U441 ( .A(n276), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U442 ( .A(n235), .B(b[7]), .ZN(n191) );
  XOR2_X1 U443 ( .A(n7), .B(n290), .Z(product[6]) );
  XNOR2_X1 U444 ( .A(n294), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U445 ( .A(n234), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U446 ( .A(n233), .B(b[3]), .ZN(n177) );
  OAI21_X1 U447 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  INV_X1 U448 ( .A(n334), .ZN(n75) );
  NOR2_X1 U449 ( .A1(n334), .A2(n44), .ZN(n39) );
  OAI22_X1 U450 ( .A1(n336), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  INV_X1 U451 ( .A(n15), .ZN(n70) );
  OAI22_X1 U452 ( .A1(n173), .A2(n343), .B1(n173), .B2(n331), .ZN(n125) );
  OAI22_X1 U453 ( .A1(n344), .A2(n174), .B1(n173), .B2(n331), .ZN(n83) );
  OAI22_X1 U454 ( .A1(n343), .A2(n175), .B1(n174), .B2(n331), .ZN(n142) );
  OAI22_X1 U455 ( .A1(n343), .A2(n176), .B1(n175), .B2(n331), .ZN(n143) );
  OAI22_X1 U456 ( .A1(n344), .A2(n177), .B1(n176), .B2(n331), .ZN(n144) );
  INV_X1 U457 ( .A(n288), .ZN(n126) );
  OAI22_X1 U458 ( .A1(n344), .A2(n179), .B1(n178), .B2(n331), .ZN(n146) );
  OAI22_X1 U459 ( .A1(n343), .A2(n178), .B1(n177), .B2(n288), .ZN(n145) );
  OAI22_X1 U460 ( .A1(n221), .A2(n229), .B1(n181), .B2(n287), .ZN(n137) );
  OAI22_X1 U461 ( .A1(n221), .A2(n180), .B1(n179), .B2(n287), .ZN(n147) );
  XNOR2_X1 U462 ( .A(n234), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U463 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U464 ( .A(n277), .B(b[1]), .ZN(n197) );
  OAI21_X1 U465 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  OAI21_X1 U466 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U467 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  XNOR2_X1 U468 ( .A(n322), .B(n1), .ZN(product[12]) );
  INV_X1 U469 ( .A(n330), .ZN(n37) );
  AOI21_X1 U470 ( .B1(n20), .B2(n339), .A(n17), .ZN(n15) );
  OAI22_X1 U471 ( .A1(n293), .A2(n193), .B1(n192), .B2(n299), .ZN(n158) );
  OAI22_X1 U472 ( .A1(n293), .A2(n195), .B1(n194), .B2(n299), .ZN(n160) );
  OAI22_X1 U473 ( .A1(n346), .A2(n194), .B1(n193), .B2(n299), .ZN(n159) );
  OAI22_X1 U474 ( .A1(n298), .A2(n196), .B1(n195), .B2(n299), .ZN(n161) );
  OAI22_X1 U475 ( .A1(n293), .A2(n231), .B1(n199), .B2(n299), .ZN(n139) );
  OAI22_X1 U476 ( .A1(n298), .A2(n197), .B1(n196), .B2(n299), .ZN(n162) );
  OAI22_X1 U477 ( .A1(n345), .A2(n192), .B1(n191), .B2(n299), .ZN(n99) );
  OAI22_X1 U478 ( .A1(n191), .A2(n346), .B1(n191), .B2(n299), .ZN(n131) );
  XNOR2_X1 U479 ( .A(n291), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U480 ( .A(n236), .B(b[6]), .ZN(n201) );
  INV_X1 U481 ( .A(n299), .ZN(n132) );
  OAI22_X1 U482 ( .A1(n223), .A2(n198), .B1(n197), .B2(n299), .ZN(n163) );
  XNOR2_X1 U483 ( .A(n291), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U484 ( .A(n236), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U485 ( .A(n289), .B(n291), .ZN(n207) );
  XNOR2_X1 U486 ( .A(n291), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U487 ( .A(n236), .B(b[3]), .ZN(n204) );
  INV_X1 U488 ( .A(n236), .ZN(n232) );
  XNOR2_X1 U489 ( .A(n236), .B(b[1]), .ZN(n206) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n74,
         n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n128,
         n129, n131, n132, n134, n135, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n229, n230, n231, n232, n233, n234, n235, n236, n244, n274,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n99), .B(n150), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n153), .B(n166), .CI(n159), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n138), .B(n155), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  CLKBUF_X2 U237 ( .A(n227), .Z(n333) );
  AND2_X1 U238 ( .A1(n118), .A2(n121), .ZN(n290) );
  BUF_X1 U239 ( .A(n227), .Z(n332) );
  NAND2_X1 U240 ( .A1(n220), .A2(n244), .ZN(n224) );
  INV_X1 U241 ( .A(n290), .ZN(n54) );
  XNOR2_X1 U242 ( .A(n234), .B(a[6]), .ZN(n274) );
  AND2_X1 U243 ( .A1(n327), .A2(n69), .ZN(product[1]) );
  XNOR2_X1 U244 ( .A(n111), .B(n276), .ZN(n104) );
  XNOR2_X1 U245 ( .A(n165), .B(n152), .ZN(n276) );
  CLKBUF_X1 U246 ( .A(n47), .Z(n277) );
  CLKBUF_X1 U247 ( .A(n45), .Z(n278) );
  CLKBUF_X1 U248 ( .A(n222), .Z(n279) );
  AOI21_X1 U249 ( .B1(n277), .B2(n39), .A(n40), .ZN(n280) );
  BUF_X2 U250 ( .A(n234), .Z(n286) );
  CLKBUF_X1 U251 ( .A(n36), .Z(n281) );
  NAND2_X1 U252 ( .A1(n111), .A2(n165), .ZN(n282) );
  NAND2_X1 U253 ( .A1(n111), .A2(n152), .ZN(n283) );
  NAND2_X1 U254 ( .A1(n165), .A2(n152), .ZN(n284) );
  NAND3_X1 U255 ( .A1(n282), .A2(n283), .A3(n284), .ZN(n103) );
  XOR2_X1 U256 ( .A(n235), .B(a[2]), .Z(n285) );
  BUF_X2 U257 ( .A(n236), .Z(n287) );
  XNOR2_X1 U258 ( .A(n104), .B(n288), .ZN(n102) );
  XNOR2_X1 U259 ( .A(n109), .B(n106), .ZN(n288) );
  AND3_X1 U260 ( .A1(n307), .A2(n306), .A3(n305), .ZN(product[15]) );
  OAI21_X1 U261 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  INV_X1 U262 ( .A(n321), .ZN(n291) );
  BUF_X1 U263 ( .A(n225), .Z(n292) );
  CLKBUF_X1 U264 ( .A(n31), .Z(n293) );
  CLKBUF_X1 U265 ( .A(n92), .Z(n294) );
  CLKBUF_X1 U266 ( .A(n70), .Z(n295) );
  NAND3_X1 U267 ( .A1(n301), .A2(n302), .A3(n303), .ZN(n296) );
  NOR2_X1 U268 ( .A1(n35), .A2(n291), .ZN(n297) );
  XNOR2_X1 U269 ( .A(n298), .B(n98), .ZN(n96) );
  XNOR2_X1 U270 ( .A(n103), .B(n105), .ZN(n298) );
  XNOR2_X1 U271 ( .A(n299), .B(n100), .ZN(n98) );
  XNOR2_X1 U272 ( .A(n145), .B(n151), .ZN(n299) );
  XOR2_X1 U273 ( .A(n85), .B(n84), .Z(n300) );
  XOR2_X1 U274 ( .A(n300), .B(n295), .Z(product[13]) );
  NAND2_X1 U275 ( .A1(n85), .A2(n84), .ZN(n301) );
  NAND2_X1 U276 ( .A1(n70), .A2(n85), .ZN(n302) );
  NAND2_X1 U277 ( .A1(n70), .A2(n84), .ZN(n303) );
  NAND3_X1 U278 ( .A1(n301), .A2(n302), .A3(n303), .ZN(n14) );
  XOR2_X1 U279 ( .A(n141), .B(n83), .Z(n304) );
  XOR2_X1 U280 ( .A(n304), .B(n296), .Z(product[14]) );
  NAND2_X1 U281 ( .A1(n141), .A2(n83), .ZN(n305) );
  NAND2_X1 U282 ( .A1(n141), .A2(n14), .ZN(n306) );
  NAND2_X1 U283 ( .A1(n83), .A2(n14), .ZN(n307) );
  NOR2_X1 U284 ( .A1(n92), .A2(n95), .ZN(n308) );
  XOR2_X1 U285 ( .A(n234), .B(a[4]), .Z(n309) );
  XNOR2_X2 U286 ( .A(n235), .B(a[4]), .ZN(n336) );
  NAND2_X1 U287 ( .A1(n145), .A2(n151), .ZN(n310) );
  NAND2_X1 U288 ( .A1(n145), .A2(n100), .ZN(n311) );
  NAND2_X1 U289 ( .A1(n151), .A2(n100), .ZN(n312) );
  NAND3_X1 U290 ( .A1(n310), .A2(n311), .A3(n312), .ZN(n97) );
  NAND2_X1 U291 ( .A1(n103), .A2(n105), .ZN(n313) );
  NAND2_X1 U292 ( .A1(n103), .A2(n98), .ZN(n314) );
  NAND2_X1 U293 ( .A1(n105), .A2(n98), .ZN(n315) );
  NAND3_X1 U294 ( .A1(n313), .A2(n314), .A3(n315), .ZN(n95) );
  CLKBUF_X1 U295 ( .A(n29), .Z(n316) );
  NAND2_X1 U296 ( .A1(n104), .A2(n109), .ZN(n317) );
  NAND2_X1 U297 ( .A1(n104), .A2(n106), .ZN(n318) );
  NAND2_X1 U298 ( .A1(n109), .A2(n106), .ZN(n319) );
  NAND3_X1 U299 ( .A1(n317), .A2(n318), .A3(n319), .ZN(n101) );
  XOR2_X1 U300 ( .A(n234), .B(a[6]), .Z(n320) );
  BUF_X2 U301 ( .A(n216), .Z(n338) );
  OR2_X1 U302 ( .A1(n294), .A2(n95), .ZN(n321) );
  AOI21_X1 U303 ( .B1(n329), .B2(n55), .A(n290), .ZN(n322) );
  NAND2_X1 U304 ( .A1(n309), .A2(n226), .ZN(n323) );
  NOR2_X1 U305 ( .A1(n102), .A2(n107), .ZN(n324) );
  NOR2_X1 U306 ( .A1(n92), .A2(n95), .ZN(n30) );
  NAND2_X1 U307 ( .A1(n285), .A2(n332), .ZN(n325) );
  NAND2_X1 U308 ( .A1(n285), .A2(n332), .ZN(n326) );
  OR2_X1 U309 ( .A1(n172), .A2(n140), .ZN(n327) );
  XNOR2_X1 U310 ( .A(n37), .B(n4), .ZN(product[9]) );
  INV_X1 U311 ( .A(n35), .ZN(n74) );
  INV_X1 U312 ( .A(n66), .ZN(n64) );
  XOR2_X1 U313 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U314 ( .A1(n328), .A2(n26), .ZN(n2) );
  INV_X1 U315 ( .A(n26), .ZN(n24) );
  AOI21_X1 U316 ( .B1(n329), .B2(n55), .A(n290), .ZN(n50) );
  NOR2_X1 U317 ( .A1(n102), .A2(n107), .ZN(n41) );
  NAND2_X1 U318 ( .A1(n331), .A2(n19), .ZN(n1) );
  XOR2_X1 U319 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U320 ( .A1(n321), .A2(n293), .ZN(n3) );
  AOI21_X1 U321 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U322 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U323 ( .A1(n76), .A2(n278), .ZN(n6) );
  INV_X1 U324 ( .A(n44), .ZN(n76) );
  XNOR2_X1 U325 ( .A(n8), .B(n55), .ZN(product[5]) );
  NAND2_X1 U326 ( .A1(n329), .A2(n54), .ZN(n8) );
  NOR2_X1 U327 ( .A1(n96), .A2(n101), .ZN(n35) );
  XNOR2_X1 U328 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U329 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U330 ( .B1(n46), .B2(n44), .A(n278), .ZN(n43) );
  XNOR2_X1 U331 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U332 ( .A1(n330), .A2(n66), .ZN(n11) );
  NAND2_X1 U333 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U334 ( .A(n48), .ZN(n77) );
  XOR2_X1 U335 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U336 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U337 ( .A(n56), .ZN(n79) );
  XOR2_X1 U338 ( .A(n10), .B(n62), .Z(product[3]) );
  INV_X1 U339 ( .A(n60), .ZN(n80) );
  INV_X1 U340 ( .A(n19), .ZN(n17) );
  OR2_X1 U341 ( .A1(n158), .A2(n146), .ZN(n105) );
  NOR2_X1 U342 ( .A1(n108), .A2(n113), .ZN(n44) );
  NOR2_X1 U343 ( .A1(n122), .A2(n123), .ZN(n56) );
  XNOR2_X1 U344 ( .A(n158), .B(n146), .ZN(n106) );
  NAND2_X1 U345 ( .A1(n108), .A2(n113), .ZN(n45) );
  NOR2_X1 U346 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U347 ( .A(n69), .ZN(n67) );
  INV_X1 U348 ( .A(n83), .ZN(n84) );
  OR2_X1 U349 ( .A1(n88), .A2(n91), .ZN(n328) );
  NAND2_X1 U350 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U351 ( .A1(n87), .A2(n86), .ZN(n19) );
  OR2_X1 U352 ( .A1(n118), .A2(n121), .ZN(n329) );
  NAND2_X1 U353 ( .A1(n114), .A2(n117), .ZN(n49) );
  OR2_X1 U354 ( .A1(n171), .A2(n164), .ZN(n330) );
  OR2_X1 U355 ( .A1(n87), .A2(n86), .ZN(n331) );
  NAND2_X1 U356 ( .A1(n122), .A2(n123), .ZN(n57) );
  AND2_X1 U357 ( .A1(n338), .A2(n132), .ZN(n164) );
  OR2_X1 U358 ( .A1(n338), .A2(n231), .ZN(n199) );
  OR2_X1 U359 ( .A1(n338), .A2(n230), .ZN(n190) );
  INV_X1 U360 ( .A(n128), .ZN(n149) );
  INV_X1 U361 ( .A(n89), .ZN(n90) );
  AND2_X1 U362 ( .A1(n338), .A2(n129), .ZN(n156) );
  INV_X1 U363 ( .A(n134), .ZN(n165) );
  AND2_X1 U364 ( .A1(n338), .A2(n320), .ZN(n148) );
  INV_X1 U365 ( .A(n125), .ZN(n141) );
  OR2_X1 U366 ( .A1(n338), .A2(n229), .ZN(n181) );
  INV_X1 U367 ( .A(n131), .ZN(n157) );
  OR2_X1 U368 ( .A1(n338), .A2(n232), .ZN(n208) );
  XNOR2_X1 U369 ( .A(n234), .B(a[6]), .ZN(n225) );
  XNOR2_X1 U370 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U371 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U372 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U373 ( .A(n233), .B(b[7]), .ZN(n173) );
  INV_X1 U374 ( .A(n135), .ZN(n244) );
  NAND2_X1 U375 ( .A1(n332), .A2(n219), .ZN(n223) );
  NAND2_X1 U376 ( .A1(n226), .A2(n218), .ZN(n222) );
  XNOR2_X1 U377 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U378 ( .A(n233), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U379 ( .A(n338), .B(n233), .ZN(n180) );
  INV_X1 U380 ( .A(n233), .ZN(n229) );
  AND2_X1 U381 ( .A1(n338), .A2(n135), .ZN(product[0]) );
  XNOR2_X1 U382 ( .A(n236), .B(a[2]), .ZN(n227) );
  NAND2_X1 U383 ( .A1(n217), .A2(n225), .ZN(n334) );
  NAND2_X1 U384 ( .A1(n217), .A2(n225), .ZN(n221) );
  CLKBUF_X1 U385 ( .A(n235), .Z(n335) );
  XNOR2_X1 U386 ( .A(n235), .B(a[4]), .ZN(n226) );
  OAI22_X1 U387 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  OAI22_X1 U388 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U389 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI22_X1 U390 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U391 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  OAI22_X1 U392 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U393 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U394 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  XOR2_X1 U395 ( .A(n233), .B(a[6]), .Z(n217) );
  INV_X1 U396 ( .A(n99), .ZN(n100) );
  INV_X1 U397 ( .A(n59), .ZN(n58) );
  AOI21_X1 U398 ( .B1(n330), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U399 ( .A(n281), .ZN(n34) );
  NAND2_X1 U400 ( .A1(n74), .A2(n281), .ZN(n4) );
  NAND2_X1 U401 ( .A1(n102), .A2(n107), .ZN(n42) );
  NOR2_X1 U402 ( .A1(n35), .A2(n308), .ZN(n28) );
  NAND2_X1 U403 ( .A1(n92), .A2(n95), .ZN(n31) );
  XNOR2_X1 U404 ( .A(n287), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U405 ( .A(n287), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U406 ( .A(n287), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U407 ( .A(n287), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U408 ( .A(n338), .B(n287), .ZN(n207) );
  XNOR2_X1 U409 ( .A(n287), .B(b[7]), .ZN(n200) );
  OAI21_X1 U410 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  NAND2_X1 U411 ( .A1(n80), .A2(n61), .ZN(n10) );
  NAND2_X1 U412 ( .A1(n124), .A2(n139), .ZN(n61) );
  NOR2_X1 U413 ( .A1(n124), .A2(n139), .ZN(n60) );
  AOI21_X1 U414 ( .B1(n29), .B2(n328), .A(n24), .ZN(n22) );
  CLKBUF_X1 U415 ( .A(n20), .Z(n337) );
  AOI21_X1 U416 ( .B1(n37), .B2(n297), .A(n316), .ZN(n27) );
  OAI22_X1 U417 ( .A1(n173), .A2(n334), .B1(n173), .B2(n274), .ZN(n125) );
  NAND2_X1 U418 ( .A1(n28), .A2(n328), .ZN(n21) );
  OAI22_X1 U419 ( .A1(n334), .A2(n174), .B1(n173), .B2(n274), .ZN(n83) );
  OAI22_X1 U420 ( .A1(n334), .A2(n175), .B1(n174), .B2(n274), .ZN(n142) );
  OAI22_X1 U421 ( .A1(n334), .A2(n176), .B1(n175), .B2(n274), .ZN(n143) );
  OAI22_X1 U422 ( .A1(n334), .A2(n177), .B1(n176), .B2(n274), .ZN(n144) );
  OAI22_X1 U423 ( .A1(n334), .A2(n179), .B1(n178), .B2(n274), .ZN(n146) );
  OAI22_X1 U424 ( .A1(n334), .A2(n178), .B1(n177), .B2(n274), .ZN(n145) );
  OAI22_X1 U425 ( .A1(n221), .A2(n229), .B1(n181), .B2(n292), .ZN(n137) );
  OAI22_X1 U426 ( .A1(n221), .A2(n180), .B1(n179), .B2(n292), .ZN(n147) );
  XOR2_X1 U427 ( .A(n236), .B(n135), .Z(n220) );
  INV_X1 U428 ( .A(n287), .ZN(n232) );
  XNOR2_X1 U429 ( .A(n287), .B(b[3]), .ZN(n204) );
  OAI21_X1 U430 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  OAI22_X1 U431 ( .A1(n182), .A2(n279), .B1(n182), .B2(n336), .ZN(n128) );
  OAI22_X1 U432 ( .A1(n323), .A2(n188), .B1(n187), .B2(n336), .ZN(n154) );
  OAI22_X1 U433 ( .A1(n279), .A2(n183), .B1(n182), .B2(n336), .ZN(n89) );
  OAI22_X1 U434 ( .A1(n222), .A2(n187), .B1(n186), .B2(n336), .ZN(n153) );
  OAI22_X1 U435 ( .A1(n323), .A2(n186), .B1(n185), .B2(n336), .ZN(n152) );
  OAI22_X1 U436 ( .A1(n222), .A2(n184), .B1(n183), .B2(n336), .ZN(n150) );
  INV_X1 U437 ( .A(n336), .ZN(n129) );
  OAI22_X1 U438 ( .A1(n323), .A2(n185), .B1(n184), .B2(n336), .ZN(n151) );
  XNOR2_X1 U439 ( .A(n235), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U440 ( .A(n235), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U441 ( .A(n235), .B(b[3]), .ZN(n195) );
  OAI22_X1 U442 ( .A1(n323), .A2(n230), .B1(n190), .B2(n336), .ZN(n138) );
  OAI22_X1 U443 ( .A1(n222), .A2(n189), .B1(n188), .B2(n336), .ZN(n155) );
  INV_X1 U444 ( .A(n335), .ZN(n231) );
  XNOR2_X1 U445 ( .A(n235), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U446 ( .A(n235), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U447 ( .A(n338), .B(n335), .ZN(n198) );
  XOR2_X1 U448 ( .A(n235), .B(a[2]), .Z(n219) );
  OAI21_X1 U449 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  NAND2_X1 U450 ( .A1(n96), .A2(n101), .ZN(n36) );
  XNOR2_X1 U451 ( .A(n235), .B(b[7]), .ZN(n191) );
  NAND2_X1 U452 ( .A1(n172), .A2(n140), .ZN(n69) );
  OAI21_X1 U453 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  AOI21_X1 U454 ( .B1(n39), .B2(n47), .A(n40), .ZN(n38) );
  INV_X1 U455 ( .A(n277), .ZN(n46) );
  OAI22_X1 U456 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  INV_X1 U457 ( .A(n324), .ZN(n75) );
  NOR2_X1 U458 ( .A1(n44), .A2(n324), .ZN(n39) );
  OAI21_X1 U459 ( .B1(n45), .B2(n41), .A(n42), .ZN(n40) );
  XNOR2_X1 U460 ( .A(n286), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U461 ( .A(b[2]), .B(n234), .ZN(n187) );
  XNOR2_X1 U462 ( .A(n286), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U463 ( .A(n286), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U464 ( .A(n234), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U465 ( .A(n286), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U466 ( .A(n338), .B(n234), .ZN(n189) );
  INV_X1 U467 ( .A(n234), .ZN(n230) );
  XOR2_X1 U468 ( .A(n234), .B(a[4]), .Z(n218) );
  XOR2_X1 U469 ( .A(n7), .B(n322), .Z(product[6]) );
  INV_X1 U470 ( .A(n15), .ZN(n70) );
  NAND2_X1 U471 ( .A1(n171), .A2(n164), .ZN(n66) );
  XNOR2_X1 U472 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U473 ( .A(n234), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U474 ( .A(n335), .B(b[1]), .ZN(n197) );
  XNOR2_X1 U475 ( .A(n287), .B(b[1]), .ZN(n206) );
  XNOR2_X1 U476 ( .A(n337), .B(n1), .ZN(product[12]) );
  INV_X1 U477 ( .A(n280), .ZN(n37) );
  AOI21_X1 U478 ( .B1(n20), .B2(n331), .A(n17), .ZN(n15) );
  OAI22_X1 U479 ( .A1(n325), .A2(n193), .B1(n192), .B2(n333), .ZN(n158) );
  OAI22_X1 U480 ( .A1(n326), .A2(n195), .B1(n194), .B2(n333), .ZN(n160) );
  OAI22_X1 U481 ( .A1(n325), .A2(n194), .B1(n193), .B2(n333), .ZN(n159) );
  OAI22_X1 U482 ( .A1(n326), .A2(n196), .B1(n195), .B2(n333), .ZN(n161) );
  OAI22_X1 U483 ( .A1(n326), .A2(n231), .B1(n199), .B2(n333), .ZN(n139) );
  OAI22_X1 U484 ( .A1(n326), .A2(n197), .B1(n196), .B2(n333), .ZN(n162) );
  OAI22_X1 U485 ( .A1(n223), .A2(n192), .B1(n191), .B2(n333), .ZN(n99) );
  OAI22_X1 U486 ( .A1(n223), .A2(n191), .B1(n191), .B2(n333), .ZN(n131) );
  INV_X1 U487 ( .A(n333), .ZN(n132) );
  OAI22_X1 U488 ( .A1(n325), .A2(n198), .B1(n197), .B2(n333), .ZN(n163) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n30, n31, n32, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n74,
         n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n131, n132, n134, n135, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n216, n217, n219, n220, n221, n222, n223, n224, n225, n227, n229,
         n230, n231, n232, n233, n234, n235, n236, n244, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n150), .B(n320), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n100), .B(n151), .CI(n145), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U110 ( .A(n153), .B(n166), .CI(n159), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n138), .B(n155), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n170), .B(n163), .CO(n123), .S(n124) );
  BUF_X1 U237 ( .A(n234), .Z(n332) );
  OR2_X1 U238 ( .A1(n172), .A2(n140), .ZN(n274) );
  XOR2_X1 U239 ( .A(n115), .B(n112), .Z(n275) );
  XOR2_X1 U240 ( .A(n110), .B(n275), .Z(n108) );
  NAND2_X1 U241 ( .A1(n110), .A2(n115), .ZN(n276) );
  NAND2_X1 U242 ( .A1(n110), .A2(n112), .ZN(n277) );
  NAND2_X1 U243 ( .A1(n115), .A2(n112), .ZN(n278) );
  NAND3_X1 U244 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n107) );
  XNOR2_X1 U245 ( .A(n104), .B(n279), .ZN(n102) );
  XNOR2_X1 U246 ( .A(n109), .B(n106), .ZN(n279) );
  XOR2_X1 U247 ( .A(n235), .B(a[4]), .Z(n280) );
  INV_X1 U248 ( .A(n34), .ZN(n281) );
  BUF_X1 U249 ( .A(n235), .Z(n288) );
  BUF_X1 U250 ( .A(n234), .Z(n333) );
  OAI21_X1 U251 ( .B1(n30), .B2(n36), .A(n31), .ZN(n282) );
  CLKBUF_X1 U252 ( .A(n326), .Z(n283) );
  NAND2_X1 U253 ( .A1(n235), .A2(n285), .ZN(n286) );
  NAND2_X1 U254 ( .A1(n284), .A2(a[2]), .ZN(n287) );
  NAND2_X1 U255 ( .A1(n286), .A2(n287), .ZN(n293) );
  INV_X1 U256 ( .A(n235), .ZN(n284) );
  INV_X1 U257 ( .A(a[2]), .ZN(n285) );
  OR2_X2 U258 ( .A1(n322), .A2(n280), .ZN(n289) );
  BUF_X2 U259 ( .A(n236), .Z(n290) );
  CLKBUF_X1 U260 ( .A(n235), .Z(n291) );
  XNOR2_X1 U261 ( .A(n158), .B(n146), .ZN(n106) );
  CLKBUF_X1 U262 ( .A(n47), .Z(n292) );
  XNOR2_X1 U263 ( .A(n236), .B(a[2]), .ZN(n294) );
  NAND2_X1 U264 ( .A1(n104), .A2(n109), .ZN(n295) );
  NAND2_X1 U265 ( .A1(n104), .A2(n106), .ZN(n296) );
  NAND2_X1 U266 ( .A1(n109), .A2(n106), .ZN(n297) );
  NAND3_X1 U267 ( .A1(n295), .A2(n296), .A3(n297), .ZN(n101) );
  CLKBUF_X1 U268 ( .A(n235), .Z(n298) );
  CLKBUF_X1 U269 ( .A(n236), .Z(n299) );
  CLKBUF_X1 U270 ( .A(n70), .Z(n300) );
  CLKBUF_X1 U271 ( .A(n40), .Z(n301) );
  BUF_X2 U272 ( .A(n227), .Z(n339) );
  XNOR2_X1 U273 ( .A(n302), .B(n308), .ZN(product[14]) );
  XNOR2_X1 U274 ( .A(n141), .B(n83), .ZN(n302) );
  AND3_X1 U275 ( .A1(n315), .A2(n314), .A3(n313), .ZN(product[15]) );
  CLKBUF_X1 U276 ( .A(n92), .Z(n304) );
  NOR2_X1 U277 ( .A1(n35), .A2(n317), .ZN(n305) );
  CLKBUF_X1 U278 ( .A(n31), .Z(n306) );
  NAND3_X1 U279 ( .A1(n312), .A2(n311), .A3(n310), .ZN(n307) );
  NAND3_X1 U280 ( .A1(n310), .A2(n311), .A3(n312), .ZN(n308) );
  XOR2_X1 U281 ( .A(n85), .B(n84), .Z(n309) );
  XOR2_X1 U282 ( .A(n309), .B(n300), .Z(product[13]) );
  NAND2_X1 U283 ( .A1(n85), .A2(n84), .ZN(n310) );
  NAND2_X1 U284 ( .A1(n70), .A2(n85), .ZN(n311) );
  NAND2_X1 U285 ( .A1(n70), .A2(n84), .ZN(n312) );
  NAND3_X1 U286 ( .A1(n310), .A2(n311), .A3(n312), .ZN(n14) );
  NAND2_X1 U287 ( .A1(n141), .A2(n83), .ZN(n313) );
  NAND2_X1 U288 ( .A1(n14), .A2(n141), .ZN(n314) );
  NAND2_X1 U289 ( .A1(n307), .A2(n83), .ZN(n315) );
  AOI21_X1 U290 ( .B1(n39), .B2(n292), .A(n301), .ZN(n316) );
  AOI21_X1 U291 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  BUF_X2 U292 ( .A(n216), .Z(n341) );
  NOR2_X1 U293 ( .A1(n92), .A2(n95), .ZN(n317) );
  NAND2_X2 U294 ( .A1(n220), .A2(n244), .ZN(n224) );
  XNOR2_X2 U295 ( .A(n235), .B(a[4]), .ZN(n340) );
  CLKBUF_X1 U296 ( .A(n282), .Z(n318) );
  CLKBUF_X1 U297 ( .A(n20), .Z(n319) );
  OAI22_X1 U298 ( .A1(n338), .A2(n192), .B1(n191), .B2(n339), .ZN(n320) );
  AOI21_X1 U299 ( .B1(n327), .B2(n55), .A(n52), .ZN(n321) );
  OR2_X2 U300 ( .A1(n322), .A2(n323), .ZN(n222) );
  XNOR2_X1 U301 ( .A(n332), .B(a[4]), .ZN(n322) );
  XOR2_X1 U302 ( .A(n235), .B(a[4]), .Z(n323) );
  OR2_X1 U303 ( .A1(n304), .A2(n95), .ZN(n324) );
  XNOR2_X1 U304 ( .A(n234), .B(a[6]), .ZN(n225) );
  NOR2_X1 U305 ( .A1(n102), .A2(n107), .ZN(n325) );
  NAND2_X1 U306 ( .A1(n217), .A2(n334), .ZN(n326) );
  INV_X1 U307 ( .A(n35), .ZN(n74) );
  XNOR2_X1 U308 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U309 ( .A1(n74), .A2(n281), .ZN(n4) );
  INV_X1 U310 ( .A(n36), .ZN(n34) );
  INV_X1 U311 ( .A(n26), .ZN(n24) );
  NAND2_X1 U312 ( .A1(n96), .A2(n101), .ZN(n36) );
  AOI21_X1 U313 ( .B1(n328), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U314 ( .A(n66), .ZN(n64) );
  NAND2_X1 U315 ( .A1(n327), .A2(n54), .ZN(n8) );
  NAND2_X1 U316 ( .A1(n330), .A2(n19), .ZN(n1) );
  XOR2_X1 U317 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U318 ( .A1(n324), .A2(n306), .ZN(n3) );
  AOI21_X1 U319 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U320 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U321 ( .A1(n76), .A2(n45), .ZN(n6) );
  INV_X1 U322 ( .A(n44), .ZN(n76) );
  XOR2_X1 U323 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U324 ( .A1(n329), .A2(n26), .ZN(n2) );
  NOR2_X1 U325 ( .A1(n96), .A2(n101), .ZN(n35) );
  XNOR2_X1 U326 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U327 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U328 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U329 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U330 ( .A1(n328), .A2(n66), .ZN(n11) );
  NAND2_X1 U331 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U332 ( .A(n48), .ZN(n77) );
  AOI21_X1 U333 ( .B1(n327), .B2(n55), .A(n52), .ZN(n50) );
  INV_X1 U334 ( .A(n54), .ZN(n52) );
  INV_X1 U335 ( .A(n19), .ZN(n17) );
  OR2_X1 U336 ( .A1(n118), .A2(n121), .ZN(n327) );
  NOR2_X1 U337 ( .A1(n108), .A2(n113), .ZN(n44) );
  NOR2_X1 U338 ( .A1(n102), .A2(n107), .ZN(n41) );
  NAND2_X1 U339 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U340 ( .A(n60), .ZN(n80) );
  INV_X1 U341 ( .A(n69), .ZN(n67) );
  OR2_X1 U342 ( .A1(n171), .A2(n164), .ZN(n328) );
  XOR2_X1 U343 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U344 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U345 ( .A(n56), .ZN(n79) );
  NAND2_X1 U346 ( .A1(n108), .A2(n113), .ZN(n45) );
  NOR2_X1 U347 ( .A1(n114), .A2(n117), .ZN(n48) );
  OR2_X1 U348 ( .A1(n88), .A2(n91), .ZN(n329) );
  NAND2_X1 U349 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U350 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U351 ( .A1(n114), .A2(n117), .ZN(n49) );
  OR2_X1 U352 ( .A1(n87), .A2(n86), .ZN(n330) );
  NAND2_X1 U353 ( .A1(n92), .A2(n95), .ZN(n31) );
  AND2_X1 U354 ( .A1(n341), .A2(n132), .ZN(n164) );
  AND2_X1 U355 ( .A1(n341), .A2(n280), .ZN(n156) );
  OAI22_X1 U356 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U357 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  OAI22_X1 U358 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  BUF_X1 U359 ( .A(n225), .Z(n335) );
  OAI22_X1 U360 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  NOR2_X1 U361 ( .A1(n122), .A2(n123), .ZN(n56) );
  NOR2_X1 U362 ( .A1(n124), .A2(n139), .ZN(n60) );
  NAND2_X1 U363 ( .A1(n122), .A2(n123), .ZN(n57) );
  AND2_X1 U364 ( .A1(n274), .A2(n69), .ZN(product[1]) );
  OR2_X1 U365 ( .A1(n341), .A2(n229), .ZN(n181) );
  OR2_X1 U366 ( .A1(n341), .A2(n231), .ZN(n199) );
  OR2_X1 U367 ( .A1(n341), .A2(n232), .ZN(n208) );
  INV_X1 U368 ( .A(n135), .ZN(n244) );
  NAND2_X1 U369 ( .A1(n217), .A2(n334), .ZN(n221) );
  AND2_X1 U370 ( .A1(n341), .A2(n135), .ZN(product[0]) );
  XNOR2_X1 U371 ( .A(n8), .B(n55), .ZN(product[5]) );
  XNOR2_X1 U372 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U373 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U374 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U375 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U376 ( .A(n341), .B(n233), .ZN(n180) );
  INV_X1 U377 ( .A(n233), .ZN(n229) );
  NAND2_X1 U378 ( .A1(n124), .A2(n139), .ZN(n61) );
  BUF_X1 U379 ( .A(n225), .Z(n334) );
  BUF_X1 U380 ( .A(n225), .Z(n336) );
  INV_X1 U381 ( .A(n134), .ZN(n165) );
  NAND2_X1 U382 ( .A1(n171), .A2(n164), .ZN(n66) );
  NAND2_X1 U383 ( .A1(n102), .A2(n107), .ZN(n42) );
  OR2_X1 U384 ( .A1(n341), .A2(n230), .ZN(n190) );
  INV_X1 U385 ( .A(n125), .ZN(n141) );
  INV_X1 U386 ( .A(n83), .ZN(n84) );
  OR2_X1 U387 ( .A1(n158), .A2(n146), .ZN(n105) );
  AND2_X1 U388 ( .A1(n341), .A2(n126), .ZN(n148) );
  INV_X1 U389 ( .A(n128), .ZN(n149) );
  INV_X1 U390 ( .A(n89), .ZN(n90) );
  OAI22_X1 U391 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  OAI22_X1 U392 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U393 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  OAI22_X1 U394 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  XOR2_X1 U395 ( .A(n233), .B(a[6]), .Z(n217) );
  NAND2_X1 U396 ( .A1(n293), .A2(n227), .ZN(n337) );
  NAND2_X1 U397 ( .A1(n219), .A2(n294), .ZN(n338) );
  NAND2_X1 U398 ( .A1(n293), .A2(n294), .ZN(n223) );
  XNOR2_X1 U399 ( .A(n236), .B(a[2]), .ZN(n227) );
  AOI21_X1 U400 ( .B1(n37), .B2(n305), .A(n318), .ZN(n27) );
  NAND2_X1 U401 ( .A1(n28), .A2(n329), .ZN(n21) );
  NOR2_X1 U402 ( .A1(n35), .A2(n317), .ZN(n28) );
  INV_X1 U403 ( .A(n99), .ZN(n100) );
  XNOR2_X1 U404 ( .A(n233), .B(b[3]), .ZN(n177) );
  XOR2_X1 U405 ( .A(n10), .B(n62), .Z(product[3]) );
  OAI21_X1 U406 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  NAND2_X1 U407 ( .A1(n172), .A2(n140), .ZN(n69) );
  INV_X1 U408 ( .A(n59), .ZN(n58) );
  NAND2_X1 U409 ( .A1(n118), .A2(n121), .ZN(n54) );
  XNOR2_X1 U410 ( .A(n233), .B(b[1]), .ZN(n179) );
  OAI21_X1 U411 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  NOR2_X1 U412 ( .A1(n92), .A2(n95), .ZN(n30) );
  INV_X1 U413 ( .A(n131), .ZN(n157) );
  XNOR2_X1 U414 ( .A(n233), .B(b[7]), .ZN(n173) );
  INV_X1 U415 ( .A(n325), .ZN(n75) );
  NOR2_X1 U416 ( .A1(n325), .A2(n44), .ZN(n39) );
  OAI21_X1 U417 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI22_X1 U418 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  AOI21_X1 U419 ( .B1(n282), .B2(n329), .A(n24), .ZN(n22) );
  OAI21_X1 U420 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  XNOR2_X1 U421 ( .A(n333), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U422 ( .A(n333), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U423 ( .A(n333), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U424 ( .A(n333), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U425 ( .A(n341), .B(n333), .ZN(n189) );
  XNOR2_X1 U426 ( .A(n333), .B(b[3]), .ZN(n186) );
  INV_X1 U427 ( .A(n332), .ZN(n230) );
  XNOR2_X1 U428 ( .A(n333), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U429 ( .A(n332), .B(b[1]), .ZN(n188) );
  XOR2_X1 U430 ( .A(n7), .B(n321), .Z(product[6]) );
  INV_X1 U431 ( .A(n292), .ZN(n46) );
  OAI21_X1 U432 ( .B1(n48), .B2(n50), .A(n49), .ZN(n47) );
  OAI22_X1 U433 ( .A1(n182), .A2(n289), .B1(n182), .B2(n340), .ZN(n128) );
  OAI22_X1 U434 ( .A1(n289), .A2(n183), .B1(n182), .B2(n340), .ZN(n89) );
  OAI22_X1 U435 ( .A1(n289), .A2(n188), .B1(n187), .B2(n340), .ZN(n154) );
  OAI22_X1 U436 ( .A1(n289), .A2(n185), .B1(n184), .B2(n340), .ZN(n151) );
  OAI22_X1 U437 ( .A1(n222), .A2(n187), .B1(n186), .B2(n340), .ZN(n153) );
  OAI22_X1 U438 ( .A1(n289), .A2(n184), .B1(n183), .B2(n340), .ZN(n150) );
  OAI22_X1 U439 ( .A1(n289), .A2(n186), .B1(n185), .B2(n340), .ZN(n152) );
  XNOR2_X1 U440 ( .A(n291), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U441 ( .A(n288), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U442 ( .A(n298), .B(b[3]), .ZN(n195) );
  OAI22_X1 U443 ( .A1(n222), .A2(n230), .B1(n190), .B2(n340), .ZN(n138) );
  OAI22_X1 U444 ( .A1(n222), .A2(n189), .B1(n188), .B2(n340), .ZN(n155) );
  XNOR2_X1 U445 ( .A(n298), .B(b[2]), .ZN(n196) );
  INV_X1 U446 ( .A(n298), .ZN(n231) );
  XNOR2_X1 U447 ( .A(n288), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U448 ( .A(n235), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U449 ( .A(n341), .B(n291), .ZN(n198) );
  XNOR2_X1 U450 ( .A(n288), .B(b[1]), .ZN(n197) );
  XOR2_X1 U451 ( .A(n235), .B(a[2]), .Z(n219) );
  INV_X1 U452 ( .A(n15), .ZN(n70) );
  OAI22_X1 U453 ( .A1(n173), .A2(n283), .B1(n173), .B2(n335), .ZN(n125) );
  OAI22_X1 U454 ( .A1(n283), .A2(n174), .B1(n173), .B2(n336), .ZN(n83) );
  OAI22_X1 U455 ( .A1(n283), .A2(n175), .B1(n174), .B2(n335), .ZN(n142) );
  OAI22_X1 U456 ( .A1(n326), .A2(n176), .B1(n175), .B2(n335), .ZN(n143) );
  OAI22_X1 U457 ( .A1(n326), .A2(n177), .B1(n176), .B2(n336), .ZN(n144) );
  OAI22_X1 U458 ( .A1(n326), .A2(n179), .B1(n178), .B2(n336), .ZN(n146) );
  OAI22_X1 U459 ( .A1(n326), .A2(n178), .B1(n177), .B2(n335), .ZN(n145) );
  INV_X1 U460 ( .A(n336), .ZN(n126) );
  OAI22_X1 U461 ( .A1(n221), .A2(n229), .B1(n181), .B2(n335), .ZN(n137) );
  OAI22_X1 U462 ( .A1(n221), .A2(n180), .B1(n179), .B2(n335), .ZN(n147) );
  XNOR2_X1 U463 ( .A(n319), .B(n1), .ZN(product[12]) );
  INV_X1 U464 ( .A(n316), .ZN(n37) );
  AOI21_X1 U465 ( .B1(n20), .B2(n330), .A(n17), .ZN(n15) );
  OAI22_X1 U466 ( .A1(n337), .A2(n193), .B1(n192), .B2(n339), .ZN(n158) );
  OAI22_X1 U467 ( .A1(n337), .A2(n195), .B1(n194), .B2(n339), .ZN(n160) );
  OAI22_X1 U468 ( .A1(n338), .A2(n194), .B1(n193), .B2(n339), .ZN(n159) );
  OAI22_X1 U469 ( .A1(n338), .A2(n196), .B1(n195), .B2(n339), .ZN(n161) );
  OAI22_X1 U470 ( .A1(n337), .A2(n231), .B1(n199), .B2(n339), .ZN(n139) );
  OAI22_X1 U471 ( .A1(n338), .A2(n197), .B1(n196), .B2(n339), .ZN(n162) );
  OAI22_X1 U472 ( .A1(n338), .A2(n192), .B1(n191), .B2(n339), .ZN(n99) );
  OAI22_X1 U473 ( .A1(n191), .A2(n337), .B1(n191), .B2(n339), .ZN(n131) );
  XNOR2_X1 U474 ( .A(n299), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U475 ( .A(n290), .B(b[6]), .ZN(n201) );
  INV_X1 U476 ( .A(n339), .ZN(n132) );
  OAI22_X1 U477 ( .A1(n223), .A2(n198), .B1(n197), .B2(n339), .ZN(n163) );
  XNOR2_X1 U478 ( .A(n299), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U479 ( .A(n290), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U480 ( .A(n341), .B(n299), .ZN(n207) );
  XNOR2_X1 U481 ( .A(n290), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U482 ( .A(n290), .B(b[3]), .ZN(n204) );
  INV_X1 U483 ( .A(n290), .ZN(n232) );
  XNOR2_X1 U484 ( .A(n290), .B(b[1]), .ZN(n206) );
  XOR2_X1 U485 ( .A(n236), .B(n135), .Z(n220) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70,
         n73, n74, n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n128, n129, n131, n132, n134, n135, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n216, n217, n218, n219, n221, n222, n223, n224, n225,
         n226, n227, n229, n230, n231, n232, n233, n234, n235, n236, n244,
         n274, n276, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n150), .B(n99), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U110 ( .A(n153), .B(n166), .CI(n159), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n160), .B(n148), .CI(n167), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  BUF_X1 U237 ( .A(n234), .Z(n301) );
  CLKBUF_X1 U238 ( .A(n55), .Z(n274) );
  AND2_X1 U239 ( .A1(n339), .A2(n69), .ZN(product[1]) );
  XNOR2_X1 U240 ( .A(n276), .B(n305), .ZN(product[14]) );
  XNOR2_X1 U241 ( .A(n141), .B(n83), .ZN(n276) );
  AND3_X1 U242 ( .A1(n312), .A2(n311), .A3(n310), .ZN(product[15]) );
  CLKBUF_X1 U243 ( .A(n236), .Z(n319) );
  CLKBUF_X2 U244 ( .A(n235), .Z(n344) );
  XNOR2_X1 U245 ( .A(n278), .B(n100), .ZN(n98) );
  XNOR2_X1 U246 ( .A(n145), .B(n151), .ZN(n278) );
  XNOR2_X1 U247 ( .A(n236), .B(a[2]), .ZN(n288) );
  NAND3_X1 U248 ( .A1(n327), .A2(n328), .A3(n329), .ZN(n279) );
  CLKBUF_X1 U249 ( .A(n36), .Z(n280) );
  CLKBUF_X1 U250 ( .A(n29), .Z(n281) );
  OR2_X2 U251 ( .A1(n282), .A2(n135), .ZN(n224) );
  XNOR2_X1 U252 ( .A(n236), .B(n135), .ZN(n282) );
  NOR2_X1 U253 ( .A1(n284), .A2(n35), .ZN(n283) );
  INV_X1 U254 ( .A(n73), .ZN(n284) );
  XNOR2_X1 U255 ( .A(n235), .B(a[4]), .ZN(n346) );
  NAND2_X1 U256 ( .A1(n70), .A2(n85), .ZN(n308) );
  NAND2_X1 U257 ( .A1(n70), .A2(n84), .ZN(n309) );
  XNOR2_X1 U258 ( .A(n110), .B(n285), .ZN(n108) );
  XNOR2_X1 U259 ( .A(n115), .B(n112), .ZN(n285) );
  INV_X1 U260 ( .A(n77), .ZN(n286) );
  XOR2_X1 U261 ( .A(a[2]), .B(n345), .Z(n287) );
  BUF_X2 U262 ( .A(n235), .Z(n345) );
  BUF_X1 U263 ( .A(n216), .Z(n289) );
  CLKBUF_X1 U264 ( .A(n221), .Z(n290) );
  NAND2_X1 U265 ( .A1(n225), .A2(n217), .ZN(n221) );
  OAI22_X1 U266 ( .A1(n221), .A2(n178), .B1(n177), .B2(n334), .ZN(n291) );
  CLKBUF_X1 U267 ( .A(n50), .Z(n292) );
  XNOR2_X1 U268 ( .A(n293), .B(n104), .ZN(n102) );
  XNOR2_X1 U269 ( .A(n109), .B(n106), .ZN(n293) );
  XNOR2_X1 U270 ( .A(n236), .B(a[2]), .ZN(n294) );
  OAI21_X1 U271 ( .B1(n286), .B2(n292), .A(n49), .ZN(n295) );
  NAND2_X1 U272 ( .A1(n233), .A2(n297), .ZN(n298) );
  NAND2_X1 U273 ( .A1(n296), .A2(a[6]), .ZN(n299) );
  NAND2_X1 U274 ( .A1(n298), .A2(n299), .ZN(n217) );
  INV_X1 U275 ( .A(n233), .ZN(n296) );
  INV_X1 U276 ( .A(a[6]), .ZN(n297) );
  CLKBUF_X1 U277 ( .A(n349), .Z(n300) );
  CLKBUF_X1 U278 ( .A(n70), .Z(n302) );
  XNOR2_X1 U279 ( .A(n303), .B(n111), .ZN(n104) );
  XNOR2_X1 U280 ( .A(n165), .B(n152), .ZN(n303) );
  NAND3_X1 U281 ( .A1(n309), .A2(n308), .A3(n307), .ZN(n304) );
  NAND3_X1 U282 ( .A1(n308), .A2(n307), .A3(n309), .ZN(n305) );
  XOR2_X1 U283 ( .A(n85), .B(n84), .Z(n306) );
  XOR2_X1 U284 ( .A(n306), .B(n302), .Z(product[13]) );
  NAND2_X1 U285 ( .A1(n85), .A2(n84), .ZN(n307) );
  NAND3_X1 U286 ( .A1(n309), .A2(n308), .A3(n307), .ZN(n14) );
  NAND2_X1 U287 ( .A1(n141), .A2(n83), .ZN(n310) );
  NAND2_X1 U288 ( .A1(n141), .A2(n14), .ZN(n311) );
  NAND2_X1 U289 ( .A1(n83), .A2(n304), .ZN(n312) );
  CLKBUF_X1 U290 ( .A(n31), .Z(n313) );
  XNOR2_X1 U291 ( .A(n314), .B(n98), .ZN(n96) );
  XNOR2_X1 U292 ( .A(n103), .B(n105), .ZN(n314) );
  NAND2_X1 U293 ( .A1(n110), .A2(n115), .ZN(n315) );
  NAND2_X1 U294 ( .A1(n110), .A2(n112), .ZN(n316) );
  NAND2_X1 U295 ( .A1(n115), .A2(n112), .ZN(n317) );
  NAND3_X1 U296 ( .A1(n315), .A2(n316), .A3(n317), .ZN(n107) );
  CLKBUF_X1 U297 ( .A(n236), .Z(n318) );
  NAND2_X1 U298 ( .A1(n291), .A2(n151), .ZN(n320) );
  NAND2_X1 U299 ( .A1(n291), .A2(n100), .ZN(n321) );
  NAND2_X1 U300 ( .A1(n151), .A2(n100), .ZN(n322) );
  NAND3_X1 U301 ( .A1(n320), .A2(n321), .A3(n322), .ZN(n97) );
  NAND2_X1 U302 ( .A1(n279), .A2(n105), .ZN(n323) );
  NAND2_X1 U303 ( .A1(n279), .A2(n98), .ZN(n324) );
  NAND2_X1 U304 ( .A1(n105), .A2(n98), .ZN(n325) );
  NAND3_X1 U305 ( .A1(n323), .A2(n324), .A3(n325), .ZN(n95) );
  NAND2_X1 U306 ( .A1(n287), .A2(n294), .ZN(n326) );
  NAND2_X1 U307 ( .A1(n165), .A2(n152), .ZN(n327) );
  NAND2_X1 U308 ( .A1(n165), .A2(n111), .ZN(n328) );
  NAND2_X1 U309 ( .A1(n152), .A2(n111), .ZN(n329) );
  NAND3_X1 U310 ( .A1(n327), .A2(n328), .A3(n329), .ZN(n103) );
  NAND2_X1 U311 ( .A1(n109), .A2(n106), .ZN(n330) );
  NAND2_X1 U312 ( .A1(n109), .A2(n104), .ZN(n331) );
  NAND2_X1 U313 ( .A1(n106), .A2(n104), .ZN(n332) );
  NAND3_X1 U314 ( .A1(n330), .A2(n331), .A3(n332), .ZN(n101) );
  INV_X1 U315 ( .A(n347), .ZN(n333) );
  INV_X2 U316 ( .A(n333), .ZN(n334) );
  CLKBUF_X1 U317 ( .A(n233), .Z(n335) );
  NOR2_X1 U318 ( .A1(n92), .A2(n95), .ZN(n336) );
  CLKBUF_X1 U319 ( .A(n20), .Z(n337) );
  AOI21_X1 U320 ( .B1(n39), .B2(n295), .A(n40), .ZN(n338) );
  XNOR2_X1 U321 ( .A(n235), .B(a[4]), .ZN(n226) );
  INV_X1 U322 ( .A(n35), .ZN(n74) );
  XNOR2_X1 U323 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U324 ( .A1(n74), .A2(n280), .ZN(n4) );
  INV_X1 U325 ( .A(n280), .ZN(n34) );
  INV_X1 U326 ( .A(n26), .ZN(n24) );
  AOI21_X1 U327 ( .B1(n341), .B2(n55), .A(n52), .ZN(n50) );
  OAI21_X1 U328 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  NAND2_X1 U329 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U330 ( .A(n60), .ZN(n80) );
  AOI21_X1 U331 ( .B1(n340), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U332 ( .A(n66), .ZN(n64) );
  NAND2_X1 U333 ( .A1(n343), .A2(n19), .ZN(n1) );
  XOR2_X1 U334 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U335 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U336 ( .A(n56), .ZN(n79) );
  XOR2_X1 U337 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U338 ( .A1(n73), .A2(n313), .ZN(n3) );
  AOI21_X1 U339 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U340 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U341 ( .A1(n76), .A2(n45), .ZN(n6) );
  INV_X1 U342 ( .A(n44), .ZN(n76) );
  XOR2_X1 U343 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U344 ( .A1(n342), .A2(n26), .ZN(n2) );
  NOR2_X1 U345 ( .A1(n336), .A2(n35), .ZN(n28) );
  XNOR2_X1 U346 ( .A(n43), .B(n5), .ZN(product[8]) );
  OAI21_X1 U347 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U348 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U349 ( .A1(n340), .A2(n66), .ZN(n11) );
  NAND2_X1 U350 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U351 ( .A(n48), .ZN(n77) );
  INV_X1 U352 ( .A(n19), .ZN(n17) );
  NOR2_X1 U353 ( .A1(n92), .A2(n95), .ZN(n30) );
  OR2_X1 U354 ( .A1(n172), .A2(n140), .ZN(n339) );
  NOR2_X1 U355 ( .A1(n108), .A2(n113), .ZN(n44) );
  XNOR2_X1 U356 ( .A(n158), .B(n146), .ZN(n106) );
  OR2_X1 U357 ( .A1(n171), .A2(n164), .ZN(n340) );
  OR2_X1 U358 ( .A1(n158), .A2(n146), .ZN(n105) );
  NAND2_X1 U359 ( .A1(n108), .A2(n113), .ZN(n45) );
  NOR2_X1 U360 ( .A1(n122), .A2(n123), .ZN(n56) );
  NOR2_X1 U361 ( .A1(n114), .A2(n117), .ZN(n48) );
  NOR2_X1 U362 ( .A1(n124), .A2(n139), .ZN(n60) );
  OR2_X1 U363 ( .A1(n118), .A2(n121), .ZN(n341) );
  INV_X1 U364 ( .A(n83), .ZN(n84) );
  OR2_X1 U365 ( .A1(n88), .A2(n91), .ZN(n342) );
  NAND2_X1 U366 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U367 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U368 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U369 ( .A1(n122), .A2(n123), .ZN(n57) );
  OR2_X1 U370 ( .A1(n87), .A2(n86), .ZN(n343) );
  AND2_X1 U371 ( .A1(n289), .A2(n132), .ZN(n164) );
  OR2_X1 U372 ( .A1(n289), .A2(n231), .ZN(n199) );
  AND2_X1 U373 ( .A1(n216), .A2(n333), .ZN(n148) );
  OR2_X1 U374 ( .A1(n289), .A2(n232), .ZN(n208) );
  INV_X1 U375 ( .A(n128), .ZN(n149) );
  INV_X1 U376 ( .A(n89), .ZN(n90) );
  AND2_X1 U377 ( .A1(n216), .A2(n129), .ZN(n156) );
  OR2_X1 U378 ( .A1(n289), .A2(n230), .ZN(n190) );
  NAND2_X1 U379 ( .A1(n219), .A2(n294), .ZN(n350) );
  INV_X1 U380 ( .A(n134), .ZN(n165) );
  INV_X1 U381 ( .A(n125), .ZN(n141) );
  OR2_X1 U382 ( .A1(n216), .A2(n229), .ZN(n181) );
  INV_X1 U383 ( .A(n135), .ZN(n244) );
  AND2_X1 U384 ( .A1(n216), .A2(n135), .ZN(product[0]) );
  INV_X1 U385 ( .A(n131), .ZN(n157) );
  NAND2_X1 U386 ( .A1(n124), .A2(n139), .ZN(n61) );
  XNOR2_X1 U387 ( .A(n236), .B(a[2]), .ZN(n227) );
  XNOR2_X1 U388 ( .A(n234), .B(a[6]), .ZN(n347) );
  XNOR2_X1 U389 ( .A(n234), .B(a[6]), .ZN(n225) );
  INV_X1 U390 ( .A(n69), .ZN(n67) );
  NAND2_X1 U391 ( .A1(n172), .A2(n140), .ZN(n69) );
  NAND2_X1 U392 ( .A1(n96), .A2(n101), .ZN(n36) );
  NOR2_X1 U393 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U394 ( .A1(n75), .A2(n42), .ZN(n5) );
  NOR2_X1 U395 ( .A1(n102), .A2(n107), .ZN(n348) );
  NOR2_X1 U396 ( .A1(n102), .A2(n107), .ZN(n41) );
  XOR2_X1 U397 ( .A(n10), .B(n62), .Z(product[3]) );
  OAI21_X1 U398 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  OAI22_X1 U399 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  NAND2_X1 U400 ( .A1(n171), .A2(n164), .ZN(n66) );
  OAI22_X1 U401 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U402 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U403 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  OAI22_X1 U404 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U405 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  NAND2_X1 U406 ( .A1(n218), .A2(n226), .ZN(n349) );
  NAND2_X1 U407 ( .A1(n218), .A2(n346), .ZN(n222) );
  XNOR2_X1 U408 ( .A(n335), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U409 ( .A(n335), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U410 ( .A(n335), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U411 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U412 ( .A(n233), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U413 ( .A(n289), .B(n233), .ZN(n180) );
  XNOR2_X1 U414 ( .A(n233), .B(b[1]), .ZN(n179) );
  INV_X1 U415 ( .A(n233), .ZN(n229) );
  NAND2_X1 U416 ( .A1(n287), .A2(n288), .ZN(n223) );
  NAND2_X1 U417 ( .A1(n341), .A2(n54), .ZN(n8) );
  INV_X1 U418 ( .A(n54), .ZN(n52) );
  OAI22_X1 U419 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U420 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  INV_X1 U421 ( .A(n59), .ZN(n58) );
  OAI21_X1 U422 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  AOI21_X1 U423 ( .B1(n37), .B2(n283), .A(n281), .ZN(n27) );
  NAND2_X1 U424 ( .A1(n28), .A2(n342), .ZN(n21) );
  INV_X1 U425 ( .A(n99), .ZN(n100) );
  XNOR2_X1 U426 ( .A(n8), .B(n274), .ZN(product[5]) );
  NAND2_X1 U427 ( .A1(n118), .A2(n121), .ZN(n54) );
  XNOR2_X1 U428 ( .A(n335), .B(b[7]), .ZN(n173) );
  AOI21_X1 U429 ( .B1(n29), .B2(n342), .A(n24), .ZN(n22) );
  OAI21_X1 U430 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  OAI22_X1 U431 ( .A1(n182), .A2(n300), .B1(n182), .B2(n226), .ZN(n128) );
  OAI22_X1 U432 ( .A1(n300), .A2(n188), .B1(n187), .B2(n346), .ZN(n154) );
  OAI22_X1 U433 ( .A1(n300), .A2(n183), .B1(n182), .B2(n226), .ZN(n89) );
  OAI22_X1 U434 ( .A1(n349), .A2(n184), .B1(n183), .B2(n346), .ZN(n150) );
  OAI22_X1 U435 ( .A1(n349), .A2(n187), .B1(n186), .B2(n346), .ZN(n153) );
  OAI22_X1 U436 ( .A1(n349), .A2(n186), .B1(n185), .B2(n346), .ZN(n152) );
  INV_X1 U437 ( .A(n226), .ZN(n129) );
  OAI22_X1 U438 ( .A1(n349), .A2(n185), .B1(n184), .B2(n226), .ZN(n151) );
  XNOR2_X1 U439 ( .A(n344), .B(b[3]), .ZN(n195) );
  OAI22_X1 U440 ( .A1(n222), .A2(n230), .B1(n190), .B2(n226), .ZN(n138) );
  OAI22_X1 U441 ( .A1(n222), .A2(n189), .B1(n188), .B2(n346), .ZN(n155) );
  XNOR2_X1 U442 ( .A(n344), .B(b[4]), .ZN(n194) );
  INV_X1 U443 ( .A(n344), .ZN(n231) );
  XNOR2_X1 U444 ( .A(n344), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U445 ( .A(n344), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U446 ( .A(n216), .B(n344), .ZN(n198) );
  XNOR2_X1 U447 ( .A(n344), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U448 ( .A(n344), .B(b[1]), .ZN(n197) );
  XNOR2_X1 U449 ( .A(n345), .B(b[7]), .ZN(n191) );
  XOR2_X1 U450 ( .A(n345), .B(a[2]), .Z(n219) );
  INV_X1 U451 ( .A(n336), .ZN(n73) );
  NAND2_X1 U452 ( .A1(n92), .A2(n95), .ZN(n31) );
  XNOR2_X1 U453 ( .A(n318), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U454 ( .A(n319), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U455 ( .A(n318), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U456 ( .A(n289), .B(n318), .ZN(n207) );
  XNOR2_X1 U457 ( .A(n319), .B(b[3]), .ZN(n204) );
  INV_X1 U458 ( .A(n319), .ZN(n232) );
  XNOR2_X1 U459 ( .A(n319), .B(b[7]), .ZN(n200) );
  INV_X1 U460 ( .A(n295), .ZN(n46) );
  AOI21_X1 U461 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U462 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  XOR2_X1 U463 ( .A(n7), .B(n292), .Z(product[6]) );
  INV_X1 U464 ( .A(n348), .ZN(n75) );
  OAI22_X1 U465 ( .A1(n173), .A2(n290), .B1(n173), .B2(n334), .ZN(n125) );
  OAI22_X1 U466 ( .A1(n290), .A2(n174), .B1(n173), .B2(n334), .ZN(n83) );
  NOR2_X1 U467 ( .A1(n348), .A2(n44), .ZN(n39) );
  OAI21_X1 U468 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  NAND2_X1 U469 ( .A1(n102), .A2(n107), .ZN(n42) );
  OAI22_X1 U470 ( .A1(n290), .A2(n175), .B1(n174), .B2(n334), .ZN(n142) );
  OAI22_X1 U471 ( .A1(n290), .A2(n176), .B1(n175), .B2(n334), .ZN(n143) );
  OAI22_X1 U472 ( .A1(n290), .A2(n177), .B1(n176), .B2(n334), .ZN(n144) );
  XNOR2_X1 U473 ( .A(n301), .B(b[7]), .ZN(n182) );
  OAI22_X1 U474 ( .A1(n221), .A2(n178), .B1(n177), .B2(n334), .ZN(n145) );
  OAI22_X1 U475 ( .A1(n221), .A2(n179), .B1(n178), .B2(n334), .ZN(n146) );
  XNOR2_X1 U476 ( .A(n234), .B(b[5]), .ZN(n184) );
  OAI22_X1 U477 ( .A1(n221), .A2(n229), .B1(n181), .B2(n347), .ZN(n137) );
  OAI22_X1 U478 ( .A1(n221), .A2(n180), .B1(n179), .B2(n347), .ZN(n147) );
  XNOR2_X1 U479 ( .A(n234), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U480 ( .A(n301), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U481 ( .A(n301), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U482 ( .A(n301), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U483 ( .A(n216), .B(n301), .ZN(n189) );
  INV_X1 U484 ( .A(n234), .ZN(n230) );
  XNOR2_X1 U485 ( .A(n234), .B(b[1]), .ZN(n188) );
  XOR2_X1 U486 ( .A(n234), .B(a[4]), .Z(n218) );
  XNOR2_X1 U487 ( .A(n319), .B(b[1]), .ZN(n206) );
  INV_X1 U488 ( .A(n15), .ZN(n70) );
  OAI22_X1 U489 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  XNOR2_X1 U490 ( .A(n318), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U491 ( .A(n337), .B(n1), .ZN(product[12]) );
  INV_X1 U492 ( .A(n338), .ZN(n37) );
  AOI21_X1 U493 ( .B1(n20), .B2(n343), .A(n17), .ZN(n15) );
  OAI22_X1 U494 ( .A1(n223), .A2(n193), .B1(n192), .B2(n227), .ZN(n158) );
  OAI22_X1 U495 ( .A1(n350), .A2(n195), .B1(n194), .B2(n227), .ZN(n160) );
  OAI22_X1 U496 ( .A1(n223), .A2(n194), .B1(n193), .B2(n294), .ZN(n159) );
  OAI22_X1 U497 ( .A1(n223), .A2(n196), .B1(n195), .B2(n227), .ZN(n161) );
  OAI22_X1 U498 ( .A1(n223), .A2(n231), .B1(n199), .B2(n227), .ZN(n139) );
  OAI22_X1 U499 ( .A1(n223), .A2(n197), .B1(n196), .B2(n288), .ZN(n162) );
  OAI22_X1 U500 ( .A1(n326), .A2(n192), .B1(n191), .B2(n227), .ZN(n99) );
  OAI22_X1 U501 ( .A1(n191), .A2(n350), .B1(n191), .B2(n227), .ZN(n131) );
  INV_X1 U502 ( .A(n288), .ZN(n132) );
  OAI22_X1 U503 ( .A1(n223), .A2(n198), .B1(n197), .B2(n227), .ZN(n163) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_10_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n56,
         n57, n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n145;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  AOI21_X1 U86 ( .B1(n33), .B2(n143), .A(n30), .ZN(n28) );
  OR2_X1 U87 ( .A1(A[0]), .A2(B[0]), .ZN(n125) );
  XOR2_X1 U88 ( .A(A[11]), .B(B[11]), .Z(n126) );
  XOR2_X1 U89 ( .A(n17), .B(n126), .Z(SUM[11]) );
  NAND2_X1 U90 ( .A1(n17), .A2(A[11]), .ZN(n127) );
  NAND2_X1 U91 ( .A1(n17), .A2(B[11]), .ZN(n128) );
  NAND2_X1 U92 ( .A1(A[11]), .A2(B[11]), .ZN(n129) );
  NAND3_X1 U93 ( .A1(n127), .A2(n128), .A3(n129), .ZN(n16) );
  INV_X1 U94 ( .A(n132), .ZN(n56) );
  CLKBUF_X1 U95 ( .A(n57), .Z(n130) );
  OR2_X2 U96 ( .A1(A[1]), .A2(B[1]), .ZN(n131) );
  AND2_X1 U97 ( .A1(A[1]), .A2(B[1]), .ZN(n132) );
  CLKBUF_X1 U98 ( .A(n49), .Z(n133) );
  AOI21_X1 U99 ( .B1(n133), .B2(n141), .A(n46), .ZN(n134) );
  CLKBUF_X1 U100 ( .A(n33), .Z(n135) );
  AOI21_X1 U101 ( .B1(n41), .B2(n142), .A(n38), .ZN(n136) );
  CLKBUF_X1 U102 ( .A(n25), .Z(n137) );
  AOI21_X1 U103 ( .B1(n131), .B2(n130), .A(n132), .ZN(n138) );
  AOI21_X1 U104 ( .B1(n131), .B2(n57), .A(n132), .ZN(n52) );
  OR2_X1 U105 ( .A1(A[3]), .A2(B[3]), .ZN(n141) );
  AOI21_X1 U106 ( .B1(n41), .B2(n142), .A(n38), .ZN(n36) );
  INV_X1 U107 ( .A(n40), .ZN(n38) );
  INV_X1 U108 ( .A(n32), .ZN(n30) );
  AOI21_X1 U109 ( .B1(n49), .B2(n141), .A(n46), .ZN(n44) );
  INV_X1 U110 ( .A(n48), .ZN(n46) );
  OAI21_X1 U111 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  NAND2_X1 U112 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U113 ( .A(n42), .ZN(n66) );
  NAND2_X1 U114 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U115 ( .A(n18), .ZN(n60) );
  OAI21_X1 U116 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  NAND2_X1 U117 ( .A1(n140), .A2(n24), .ZN(n3) );
  NAND2_X1 U118 ( .A1(n141), .A2(n48), .ZN(n9) );
  NAND2_X1 U119 ( .A1(n142), .A2(n40), .ZN(n7) );
  XOR2_X1 U120 ( .A(n138), .B(n10), .Z(SUM[2]) );
  NAND2_X1 U121 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U122 ( .A(n50), .ZN(n68) );
  XOR2_X1 U123 ( .A(n28), .B(n4), .Z(SUM[8]) );
  NAND2_X1 U124 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U125 ( .A(n26), .ZN(n62) );
  XOR2_X1 U126 ( .A(n136), .B(n6), .Z(SUM[6]) );
  NAND2_X1 U127 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U128 ( .A(n34), .ZN(n64) );
  XNOR2_X1 U129 ( .A(n135), .B(n5), .ZN(SUM[7]) );
  NAND2_X1 U130 ( .A1(n143), .A2(n32), .ZN(n5) );
  INV_X1 U131 ( .A(n59), .ZN(n57) );
  XNOR2_X1 U132 ( .A(n11), .B(n130), .ZN(SUM[1]) );
  NAND2_X1 U133 ( .A1(n131), .A2(n56), .ZN(n11) );
  INV_X1 U134 ( .A(n24), .ZN(n22) );
  XNOR2_X1 U135 ( .A(n13), .B(n139), .ZN(SUM[15]) );
  XNOR2_X1 U136 ( .A(B[15]), .B(A[15]), .ZN(n139) );
  NOR2_X1 U137 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U138 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  OR2_X1 U139 ( .A1(A[9]), .A2(B[9]), .ZN(n140) );
  OR2_X1 U140 ( .A1(A[5]), .A2(B[5]), .ZN(n142) );
  NOR2_X1 U141 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U142 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U144 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U145 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U146 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U147 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U148 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  NAND2_X1 U149 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  OR2_X1 U150 ( .A1(A[7]), .A2(B[7]), .ZN(n143) );
  NAND2_X1 U151 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U152 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U153 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  AND2_X1 U154 ( .A1(n125), .A2(n59), .ZN(SUM[0]) );
  AOI21_X1 U155 ( .B1(n137), .B2(n140), .A(n22), .ZN(n145) );
  XNOR2_X1 U156 ( .A(n137), .B(n3), .ZN(SUM[9]) );
  XNOR2_X1 U157 ( .A(n41), .B(n7), .ZN(SUM[5]) );
  AOI21_X1 U158 ( .B1(n25), .B2(n140), .A(n22), .ZN(n20) );
  OAI21_X1 U159 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  XOR2_X1 U160 ( .A(n134), .B(n8), .Z(SUM[4]) );
  XNOR2_X1 U161 ( .A(n133), .B(n9), .ZN(SUM[3]) );
  XOR2_X1 U162 ( .A(n145), .B(n2), .Z(SUM[10]) );
  NAND2_X1 U163 ( .A1(A[0]), .A2(B[0]), .ZN(n59) );
  OAI21_X1 U164 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X1 U165 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
endmodule


module add_layer_WIDTH16_10 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_10_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_9_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n56,
         n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  AND2_X1 U86 ( .A1(A[1]), .A2(B[1]), .ZN(n132) );
  AOI21_X1 U87 ( .B1(n41), .B2(n141), .A(n38), .ZN(n36) );
  INV_X1 U88 ( .A(n132), .ZN(n56) );
  OR2_X1 U89 ( .A1(A[0]), .A2(B[0]), .ZN(n125) );
  XOR2_X1 U90 ( .A(A[11]), .B(B[11]), .Z(n126) );
  XOR2_X1 U91 ( .A(n17), .B(n126), .Z(SUM[11]) );
  NAND2_X1 U92 ( .A1(n17), .A2(A[11]), .ZN(n127) );
  NAND2_X1 U93 ( .A1(n17), .A2(B[11]), .ZN(n128) );
  NAND2_X1 U94 ( .A1(A[11]), .A2(B[11]), .ZN(n129) );
  NAND3_X1 U95 ( .A1(n127), .A2(n128), .A3(n129), .ZN(n16) );
  OR2_X2 U96 ( .A1(A[1]), .A2(B[1]), .ZN(n139) );
  AOI21_X1 U97 ( .B1(n139), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U98 ( .B1(n139), .B2(n131), .A(n132), .ZN(n52) );
  AND2_X1 U99 ( .A1(A[0]), .A2(B[0]), .ZN(n131) );
  CLKBUF_X1 U100 ( .A(n49), .Z(n133) );
  CLKBUF_X1 U101 ( .A(n33), .Z(n134) );
  CLKBUF_X1 U102 ( .A(n25), .Z(n135) );
  AOI21_X1 U103 ( .B1(n133), .B2(n142), .A(n46), .ZN(n136) );
  AOI21_X1 U104 ( .B1(n135), .B2(n143), .A(n22), .ZN(n137) );
  AOI21_X1 U105 ( .B1(n134), .B2(n144), .A(n30), .ZN(n138) );
  INV_X1 U106 ( .A(n24), .ZN(n22) );
  INV_X1 U107 ( .A(n48), .ZN(n46) );
  INV_X1 U108 ( .A(n40), .ZN(n38) );
  AOI21_X1 U109 ( .B1(n33), .B2(n144), .A(n30), .ZN(n28) );
  INV_X1 U110 ( .A(n32), .ZN(n30) );
  NAND2_X1 U111 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U112 ( .A(n42), .ZN(n66) );
  NAND2_X1 U113 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U114 ( .A(n34), .ZN(n64) );
  NAND2_X1 U115 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U116 ( .A(n26), .ZN(n62) );
  NAND2_X1 U117 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U118 ( .A(n18), .ZN(n60) );
  NAND2_X1 U119 ( .A1(n141), .A2(n40), .ZN(n7) );
  NAND2_X1 U120 ( .A1(n142), .A2(n48), .ZN(n9) );
  NAND2_X1 U121 ( .A1(n143), .A2(n24), .ZN(n3) );
  XNOR2_X1 U122 ( .A(n134), .B(n5), .ZN(SUM[7]) );
  NAND2_X1 U123 ( .A1(n144), .A2(n32), .ZN(n5) );
  XNOR2_X1 U124 ( .A(n11), .B(n131), .ZN(SUM[1]) );
  NAND2_X1 U125 ( .A1(n139), .A2(n56), .ZN(n11) );
  NAND2_X1 U126 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U127 ( .A(n50), .ZN(n68) );
  XNOR2_X1 U128 ( .A(n13), .B(n140), .ZN(SUM[15]) );
  XNOR2_X1 U129 ( .A(B[15]), .B(A[15]), .ZN(n140) );
  NOR2_X1 U130 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  NOR2_X1 U131 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U132 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U133 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U134 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U135 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U136 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U137 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U138 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  OR2_X1 U139 ( .A1(A[5]), .A2(B[5]), .ZN(n141) );
  OR2_X1 U140 ( .A1(A[3]), .A2(B[3]), .ZN(n142) );
  OR2_X1 U141 ( .A1(A[9]), .A2(B[9]), .ZN(n143) );
  OR2_X1 U142 ( .A1(A[7]), .A2(B[7]), .ZN(n144) );
  NAND2_X1 U143 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  NAND2_X1 U144 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U145 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U146 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U147 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  AND2_X1 U148 ( .A1(n125), .A2(n59), .ZN(SUM[0]) );
  XOR2_X1 U149 ( .A(n36), .B(n6), .Z(SUM[6]) );
  OAI21_X1 U150 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U151 ( .A(n41), .B(n7), .ZN(SUM[5]) );
  XOR2_X1 U152 ( .A(n136), .B(n8), .Z(SUM[4]) );
  OAI21_X1 U153 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  AOI21_X1 U154 ( .B1(n49), .B2(n142), .A(n46), .ZN(n44) );
  XNOR2_X1 U155 ( .A(n133), .B(n9), .ZN(SUM[3]) );
  NAND2_X1 U156 ( .A1(A[0]), .A2(B[0]), .ZN(n59) );
  XNOR2_X1 U157 ( .A(n135), .B(n3), .ZN(SUM[9]) );
  XOR2_X1 U158 ( .A(n130), .B(n10), .Z(SUM[2]) );
  XOR2_X1 U159 ( .A(n137), .B(n2), .Z(SUM[10]) );
  AOI21_X1 U160 ( .B1(n25), .B2(n143), .A(n22), .ZN(n20) );
  OAI21_X1 U161 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X1 U162 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U163 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U164 ( .A(n138), .B(n4), .Z(SUM[8]) );
endmodule


module add_layer_WIDTH16_9 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_9_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n16, n21, n22,
         n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37, n38, n39, n40,
         n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55, n56, n57, n61,
         n64, n65, n67, n69, n71, n73, n75, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n160,
         n161, n162;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n15), .CO(n14), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n16), .CO(n15), .S(SUM[13]) );
  OR2_X1 U94 ( .A1(A[0]), .A2(B[0]), .ZN(n132) );
  CLKBUF_X1 U95 ( .A(n65), .Z(n133) );
  XOR2_X1 U96 ( .A(A[12]), .B(B[12]), .Z(n134) );
  XOR2_X1 U97 ( .A(n133), .B(n134), .Z(SUM[12]) );
  NAND2_X1 U98 ( .A1(n65), .A2(A[12]), .ZN(n135) );
  NAND2_X1 U99 ( .A1(n65), .A2(B[12]), .ZN(n136) );
  NAND2_X1 U100 ( .A1(A[12]), .A2(B[12]), .ZN(n137) );
  NAND3_X1 U101 ( .A1(n136), .A2(n135), .A3(n137), .ZN(n16) );
  OAI21_X1 U102 ( .B1(n139), .B2(n138), .A(n21), .ZN(n65) );
  INV_X1 U103 ( .A(n162), .ZN(n138) );
  INV_X1 U104 ( .A(n22), .ZN(n139) );
  OR2_X1 U105 ( .A1(A[1]), .A2(B[1]), .ZN(n140) );
  INV_X1 U106 ( .A(n61), .ZN(n141) );
  INV_X1 U107 ( .A(n143), .ZN(n61) );
  AND2_X1 U108 ( .A1(A[1]), .A2(B[1]), .ZN(n143) );
  AND2_X1 U109 ( .A1(A[0]), .A2(B[0]), .ZN(n142) );
  CLKBUF_X1 U110 ( .A(n30), .Z(n144) );
  CLKBUF_X1 U111 ( .A(n46), .Z(n145) );
  CLKBUF_X1 U112 ( .A(n54), .Z(n146) );
  AOI21_X1 U113 ( .B1(n144), .B2(n160), .A(n27), .ZN(n147) );
  CLKBUF_X1 U114 ( .A(n38), .Z(n148) );
  AOI21_X1 U115 ( .B1(n146), .B2(n157), .A(n51), .ZN(n149) );
  AOI21_X1 U116 ( .B1(n145), .B2(n155), .A(n43), .ZN(n150) );
  CLKBUF_X1 U117 ( .A(n22), .Z(n151) );
  AOI21_X1 U118 ( .B1(n54), .B2(n157), .A(n51), .ZN(n49) );
  AOI21_X1 U119 ( .B1(n46), .B2(n155), .A(n43), .ZN(n41) );
  AOI21_X1 U120 ( .B1(n38), .B2(n161), .A(n35), .ZN(n152) );
  AOI21_X1 U121 ( .B1(n158), .B2(n142), .A(n143), .ZN(n153) );
  XNOR2_X1 U122 ( .A(n154), .B(n142), .ZN(SUM[1]) );
  NAND2_X1 U123 ( .A1(n140), .A2(n61), .ZN(n154) );
  OR2_X1 U124 ( .A1(A[5]), .A2(B[5]), .ZN(n155) );
  INV_X1 U125 ( .A(n29), .ZN(n27) );
  INV_X1 U126 ( .A(n37), .ZN(n35) );
  INV_X1 U127 ( .A(n45), .ZN(n43) );
  INV_X1 U128 ( .A(n53), .ZN(n51) );
  AOI21_X1 U129 ( .B1(n140), .B2(n142), .A(n141), .ZN(n57) );
  NAND2_X1 U130 ( .A1(n67), .A2(n24), .ZN(n3) );
  INV_X1 U131 ( .A(n23), .ZN(n67) );
  NAND2_X1 U132 ( .A1(n73), .A2(n48), .ZN(n9) );
  INV_X1 U133 ( .A(n47), .ZN(n73) );
  NAND2_X1 U134 ( .A1(n69), .A2(n32), .ZN(n5) );
  INV_X1 U135 ( .A(n31), .ZN(n69) );
  NAND2_X1 U136 ( .A1(n162), .A2(n21), .ZN(n2) );
  NAND2_X1 U137 ( .A1(n161), .A2(n37), .ZN(n6) );
  NAND2_X1 U138 ( .A1(n157), .A2(n53), .ZN(n10) );
  NAND2_X1 U139 ( .A1(n155), .A2(n45), .ZN(n8) );
  NAND2_X1 U140 ( .A1(n160), .A2(n29), .ZN(n4) );
  NAND2_X1 U141 ( .A1(n71), .A2(n40), .ZN(n7) );
  INV_X1 U142 ( .A(n39), .ZN(n71) );
  NAND2_X1 U143 ( .A1(n75), .A2(n56), .ZN(n11) );
  INV_X1 U144 ( .A(n55), .ZN(n75) );
  XNOR2_X1 U145 ( .A(n14), .B(n156), .ZN(SUM[15]) );
  XNOR2_X1 U146 ( .A(B[15]), .B(A[15]), .ZN(n156) );
  OR2_X1 U147 ( .A1(A[3]), .A2(B[3]), .ZN(n157) );
  NOR2_X1 U148 ( .A1(A[6]), .A2(B[6]), .ZN(n39) );
  NOR2_X1 U149 ( .A1(A[8]), .A2(B[8]), .ZN(n31) );
  NOR2_X1 U150 ( .A1(A[2]), .A2(B[2]), .ZN(n55) );
  NOR2_X1 U151 ( .A1(A[4]), .A2(B[4]), .ZN(n47) );
  NOR2_X1 U152 ( .A1(A[10]), .A2(B[10]), .ZN(n23) );
  OR2_X1 U153 ( .A1(A[1]), .A2(B[1]), .ZN(n158) );
  AND2_X1 U154 ( .A1(n132), .A2(n64), .ZN(SUM[0]) );
  NAND2_X1 U155 ( .A1(A[9]), .A2(B[9]), .ZN(n29) );
  NAND2_X1 U156 ( .A1(A[7]), .A2(B[7]), .ZN(n37) );
  NAND2_X1 U157 ( .A1(A[5]), .A2(B[5]), .ZN(n45) );
  NAND2_X1 U158 ( .A1(A[3]), .A2(B[3]), .ZN(n53) );
  NAND2_X1 U159 ( .A1(A[11]), .A2(B[11]), .ZN(n21) );
  OR2_X1 U160 ( .A1(A[9]), .A2(B[9]), .ZN(n160) );
  OR2_X1 U161 ( .A1(A[7]), .A2(B[7]), .ZN(n161) );
  OR2_X1 U162 ( .A1(A[11]), .A2(B[11]), .ZN(n162) );
  NAND2_X1 U163 ( .A1(A[6]), .A2(B[6]), .ZN(n40) );
  NAND2_X1 U164 ( .A1(A[8]), .A2(B[8]), .ZN(n32) );
  NAND2_X1 U165 ( .A1(A[2]), .A2(B[2]), .ZN(n56) );
  NAND2_X1 U166 ( .A1(A[4]), .A2(B[4]), .ZN(n48) );
  NAND2_X1 U167 ( .A1(A[10]), .A2(B[10]), .ZN(n24) );
  XOR2_X1 U168 ( .A(n150), .B(n7), .Z(SUM[6]) );
  XOR2_X1 U169 ( .A(n33), .B(n5), .Z(SUM[8]) );
  AOI21_X1 U170 ( .B1(n148), .B2(n161), .A(n35), .ZN(n33) );
  XNOR2_X1 U171 ( .A(n145), .B(n8), .ZN(SUM[5]) );
  XNOR2_X1 U172 ( .A(n148), .B(n6), .ZN(SUM[7]) );
  NAND2_X1 U173 ( .A1(A[0]), .A2(B[0]), .ZN(n64) );
  OAI21_X1 U174 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U175 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  XOR2_X1 U176 ( .A(n149), .B(n9), .Z(SUM[4]) );
  XNOR2_X1 U177 ( .A(n144), .B(n4), .ZN(SUM[9]) );
  XNOR2_X1 U178 ( .A(n146), .B(n10), .ZN(SUM[3]) );
  OAI21_X1 U179 ( .B1(n152), .B2(n31), .A(n32), .ZN(n30) );
  OAI21_X1 U180 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
  XOR2_X1 U181 ( .A(n147), .B(n3), .Z(SUM[10]) );
  XNOR2_X1 U182 ( .A(n151), .B(n2), .ZN(SUM[11]) );
  AOI21_X1 U183 ( .B1(n30), .B2(n160), .A(n27), .ZN(n25) );
  OAI21_X1 U184 ( .B1(n153), .B2(n55), .A(n56), .ZN(n54) );
  XOR2_X1 U185 ( .A(n57), .B(n11), .Z(SUM[2]) );
endmodule


module add_layer_WIDTH16_3 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_3_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_3 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_3 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_3 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_10 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_9 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_3 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_3 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12 \genblk1[0].mult  ( .clk(clk), 
        .ia({\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11 \genblk1[1].mult  ( .clk(clk), 
        .ia({\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10 \genblk1[2].mult  ( .clk(clk), 
        .ia({\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9 \genblk1[3].mult  ( .clk(clk), .ia(
        {\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_3 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n31, n32, n34, n35, n36, n37, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n73, n74,
         n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n129, n131, n132, n134, n135, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n216, n217, n218, n219, n221, n222, n223, n224, n225, n226,
         n227, n229, n230, n231, n232, n233, n234, n235, n236, n244, n274,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n157), .B(n99), .CI(n150), .CO(n93), .S(n94) );
  FA_X1 U103 ( .A(n145), .B(n151), .CI(n100), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U110 ( .A(n159), .B(n166), .CI(n153), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  CLKBUF_X3 U237 ( .A(n226), .Z(n319) );
  CLKBUF_X1 U238 ( .A(n47), .Z(n274) );
  BUF_X2 U239 ( .A(n227), .Z(n327) );
  OR2_X1 U240 ( .A1(n88), .A2(n91), .ZN(n323) );
  AND2_X1 U241 ( .A1(n322), .A2(n69), .ZN(product[1]) );
  INV_X1 U242 ( .A(n281), .ZN(n276) );
  INV_X1 U243 ( .A(n281), .ZN(n282) );
  XOR2_X1 U244 ( .A(n233), .B(a[6]), .Z(n277) );
  BUF_X2 U245 ( .A(n234), .Z(n278) );
  NAND2_X1 U246 ( .A1(n217), .A2(n225), .ZN(n221) );
  OR2_X2 U247 ( .A1(n279), .A2(n135), .ZN(n224) );
  XNOR2_X1 U248 ( .A(n236), .B(n135), .ZN(n279) );
  INV_X1 U249 ( .A(n135), .ZN(n244) );
  BUF_X1 U250 ( .A(n218), .Z(n280) );
  INV_X1 U251 ( .A(n235), .ZN(n281) );
  XNOR2_X1 U252 ( .A(n235), .B(a[4]), .ZN(n283) );
  XNOR2_X1 U253 ( .A(n284), .B(n306), .ZN(product[14]) );
  XNOR2_X1 U254 ( .A(n141), .B(n83), .ZN(n284) );
  AND3_X1 U255 ( .A1(n314), .A2(n313), .A3(n312), .ZN(product[15]) );
  XNOR2_X1 U256 ( .A(n104), .B(n286), .ZN(n102) );
  XNOR2_X1 U257 ( .A(n109), .B(n106), .ZN(n286) );
  XNOR2_X1 U258 ( .A(n287), .B(n98), .ZN(n96) );
  XNOR2_X1 U259 ( .A(n103), .B(n105), .ZN(n287) );
  OAI21_X2 U260 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  BUF_X1 U261 ( .A(n236), .Z(n288) );
  CLKBUF_X1 U262 ( .A(n236), .Z(n289) );
  NAND2_X1 U263 ( .A1(n98), .A2(n103), .ZN(n290) );
  NAND2_X1 U264 ( .A1(n98), .A2(n105), .ZN(n291) );
  NAND2_X1 U265 ( .A1(n103), .A2(n105), .ZN(n292) );
  NAND3_X1 U266 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n95) );
  NAND2_X1 U267 ( .A1(n104), .A2(n109), .ZN(n293) );
  NAND2_X1 U268 ( .A1(n104), .A2(n106), .ZN(n294) );
  NAND2_X1 U269 ( .A1(n109), .A2(n106), .ZN(n295) );
  NAND3_X1 U270 ( .A1(n293), .A2(n294), .A3(n295), .ZN(n101) );
  XOR2_X1 U271 ( .A(n115), .B(n112), .Z(n296) );
  XOR2_X1 U272 ( .A(n110), .B(n296), .Z(n108) );
  NAND2_X1 U273 ( .A1(n110), .A2(n115), .ZN(n297) );
  NAND2_X1 U274 ( .A1(n110), .A2(n112), .ZN(n298) );
  NAND2_X1 U275 ( .A1(n115), .A2(n112), .ZN(n299) );
  NAND3_X1 U276 ( .A1(n297), .A2(n298), .A3(n299), .ZN(n107) );
  CLKBUF_X1 U277 ( .A(n36), .Z(n300) );
  CLKBUF_X1 U278 ( .A(n315), .Z(n301) );
  CLKBUF_X1 U279 ( .A(n70), .Z(n302) );
  NOR2_X1 U280 ( .A1(n35), .A2(n317), .ZN(n303) );
  XNOR2_X1 U281 ( .A(n234), .B(a[6]), .ZN(n304) );
  BUF_X2 U282 ( .A(n225), .Z(n330) );
  NAND3_X1 U283 ( .A1(n311), .A2(n310), .A3(n309), .ZN(n305) );
  NAND3_X1 U284 ( .A1(n311), .A2(n310), .A3(n309), .ZN(n306) );
  CLKBUF_X1 U285 ( .A(n20), .Z(n307) );
  XOR2_X1 U286 ( .A(n85), .B(n84), .Z(n308) );
  XOR2_X1 U287 ( .A(n308), .B(n302), .Z(product[13]) );
  NAND2_X1 U288 ( .A1(n85), .A2(n84), .ZN(n309) );
  NAND2_X1 U289 ( .A1(n70), .A2(n85), .ZN(n310) );
  NAND2_X1 U290 ( .A1(n70), .A2(n84), .ZN(n311) );
  NAND3_X1 U291 ( .A1(n310), .A2(n309), .A3(n311), .ZN(n14) );
  NAND2_X1 U292 ( .A1(n141), .A2(n83), .ZN(n312) );
  NAND2_X1 U293 ( .A1(n14), .A2(n141), .ZN(n313) );
  NAND2_X1 U294 ( .A1(n83), .A2(n305), .ZN(n314) );
  AOI21_X1 U295 ( .B1(n47), .B2(n39), .A(n40), .ZN(n315) );
  NOR2_X1 U296 ( .A1(n92), .A2(n95), .ZN(n316) );
  NOR2_X1 U297 ( .A1(n92), .A2(n95), .ZN(n317) );
  AOI21_X1 U298 ( .B1(n326), .B2(n55), .A(n52), .ZN(n318) );
  XNOR2_X1 U299 ( .A(n235), .B(a[4]), .ZN(n226) );
  BUF_X2 U300 ( .A(n216), .Z(n334) );
  NOR2_X1 U301 ( .A1(n102), .A2(n107), .ZN(n320) );
  XOR2_X1 U302 ( .A(n43), .B(n321), .Z(product[8]) );
  AND2_X1 U303 ( .A1(n75), .A2(n42), .ZN(n321) );
  NOR2_X1 U304 ( .A1(n108), .A2(n113), .ZN(n44) );
  OR2_X1 U305 ( .A1(n172), .A2(n140), .ZN(n322) );
  INV_X1 U306 ( .A(n35), .ZN(n74) );
  XNOR2_X1 U307 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U308 ( .A1(n74), .A2(n300), .ZN(n4) );
  INV_X1 U309 ( .A(n300), .ZN(n34) );
  INV_X1 U310 ( .A(n66), .ZN(n64) );
  INV_X1 U311 ( .A(n26), .ZN(n24) );
  NOR2_X1 U312 ( .A1(n102), .A2(n107), .ZN(n41) );
  NOR2_X1 U313 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U314 ( .A1(n325), .A2(n19), .ZN(n1) );
  XOR2_X1 U315 ( .A(n46), .B(n6), .Z(product[7]) );
  INV_X1 U316 ( .A(n44), .ZN(n76) );
  XOR2_X1 U317 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U318 ( .A1(n73), .A2(n31), .ZN(n3) );
  AOI21_X1 U319 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U320 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U321 ( .A1(n323), .A2(n26), .ZN(n2) );
  XNOR2_X1 U322 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U323 ( .A1(n324), .A2(n66), .ZN(n11) );
  NAND2_X1 U324 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U325 ( .A(n48), .ZN(n77) );
  INV_X1 U326 ( .A(n19), .ZN(n17) );
  XNOR2_X1 U327 ( .A(n158), .B(n146), .ZN(n106) );
  OR2_X1 U328 ( .A1(n158), .A2(n146), .ZN(n105) );
  XOR2_X1 U329 ( .A(n10), .B(n62), .Z(product[3]) );
  INV_X1 U330 ( .A(n60), .ZN(n80) );
  XOR2_X1 U331 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U332 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U333 ( .A(n56), .ZN(n79) );
  NAND2_X1 U334 ( .A1(n172), .A2(n140), .ZN(n69) );
  NOR2_X1 U335 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U336 ( .A(n83), .ZN(n84) );
  NAND2_X1 U337 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U338 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U339 ( .A1(n114), .A2(n117), .ZN(n49) );
  OR2_X1 U340 ( .A1(n171), .A2(n164), .ZN(n324) );
  OR2_X1 U341 ( .A1(n87), .A2(n86), .ZN(n325) );
  OR2_X1 U342 ( .A1(n118), .A2(n121), .ZN(n326) );
  AND2_X1 U343 ( .A1(n334), .A2(n132), .ZN(n164) );
  OR2_X1 U344 ( .A1(n334), .A2(n232), .ZN(n208) );
  OAI22_X1 U345 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  INV_X1 U346 ( .A(n128), .ZN(n149) );
  INV_X1 U347 ( .A(n89), .ZN(n90) );
  AND2_X1 U348 ( .A1(n334), .A2(n129), .ZN(n156) );
  OAI22_X1 U349 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OR2_X1 U350 ( .A1(n334), .A2(n230), .ZN(n190) );
  OAI22_X1 U351 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  NOR2_X1 U352 ( .A1(n124), .A2(n139), .ZN(n60) );
  NOR2_X1 U353 ( .A1(n122), .A2(n123), .ZN(n56) );
  NAND2_X1 U354 ( .A1(n124), .A2(n139), .ZN(n61) );
  INV_X1 U355 ( .A(n131), .ZN(n157) );
  AND2_X1 U356 ( .A1(n334), .A2(n126), .ZN(n148) );
  INV_X1 U357 ( .A(n125), .ZN(n141) );
  NAND2_X1 U358 ( .A1(n122), .A2(n123), .ZN(n57) );
  INV_X1 U359 ( .A(n99), .ZN(n100) );
  OR2_X1 U360 ( .A1(n334), .A2(n229), .ZN(n181) );
  OR2_X1 U361 ( .A1(n334), .A2(n231), .ZN(n199) );
  XNOR2_X1 U362 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U363 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U364 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U365 ( .A(n334), .B(n233), .ZN(n180) );
  INV_X1 U366 ( .A(n233), .ZN(n229) );
  AND2_X1 U367 ( .A1(n334), .A2(n135), .ZN(product[0]) );
  XNOR2_X1 U368 ( .A(n236), .B(a[2]), .ZN(n227) );
  NAND2_X1 U369 ( .A1(n280), .A2(n319), .ZN(n333) );
  NAND2_X1 U370 ( .A1(n280), .A2(n319), .ZN(n332) );
  NAND2_X1 U371 ( .A1(n218), .A2(n283), .ZN(n222) );
  OAI21_X1 U372 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  NAND2_X1 U373 ( .A1(n76), .A2(n45), .ZN(n6) );
  XNOR2_X1 U374 ( .A(n233), .B(b[6]), .ZN(n174) );
  OAI22_X1 U375 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U376 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  NAND2_X1 U377 ( .A1(n326), .A2(n54), .ZN(n8) );
  INV_X1 U378 ( .A(n54), .ZN(n52) );
  NAND2_X1 U379 ( .A1(n277), .A2(n330), .ZN(n328) );
  NAND2_X1 U380 ( .A1(n277), .A2(n304), .ZN(n329) );
  XOR2_X1 U381 ( .A(n233), .B(a[6]), .Z(n217) );
  XNOR2_X1 U382 ( .A(n234), .B(a[6]), .ZN(n225) );
  NAND2_X1 U383 ( .A1(n108), .A2(n113), .ZN(n45) );
  NAND2_X1 U384 ( .A1(n80), .A2(n61), .ZN(n10) );
  OAI21_X1 U385 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  NAND2_X1 U386 ( .A1(n227), .A2(n219), .ZN(n331) );
  NAND2_X1 U387 ( .A1(n219), .A2(n227), .ZN(n223) );
  NAND2_X1 U388 ( .A1(n28), .A2(n323), .ZN(n21) );
  OAI21_X1 U389 ( .B1(n316), .B2(n36), .A(n31), .ZN(n29) );
  NOR2_X1 U390 ( .A1(n317), .A2(n35), .ZN(n28) );
  XNOR2_X1 U391 ( .A(n233), .B(b[7]), .ZN(n173) );
  XNOR2_X1 U392 ( .A(n8), .B(n55), .ZN(product[5]) );
  INV_X1 U393 ( .A(n134), .ZN(n165) );
  OAI22_X1 U394 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  AOI21_X1 U395 ( .B1(n324), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U396 ( .A(n69), .ZN(n67) );
  INV_X1 U397 ( .A(n59), .ZN(n58) );
  OAI22_X1 U398 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  XOR2_X1 U399 ( .A(n235), .B(a[2]), .Z(n219) );
  INV_X1 U400 ( .A(n276), .ZN(n231) );
  XNOR2_X1 U401 ( .A(n235), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U402 ( .A(n282), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U403 ( .A(n276), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U404 ( .A(n282), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U405 ( .A(n276), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U406 ( .A(n334), .B(n276), .ZN(n198) );
  NAND2_X1 U407 ( .A1(n118), .A2(n121), .ZN(n54) );
  OAI22_X1 U408 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  AOI21_X1 U409 ( .B1(n37), .B2(n303), .A(n29), .ZN(n27) );
  OAI22_X1 U410 ( .A1(n173), .A2(n328), .B1(n173), .B2(n330), .ZN(n125) );
  OAI22_X1 U411 ( .A1(n329), .A2(n174), .B1(n173), .B2(n304), .ZN(n83) );
  AOI21_X1 U412 ( .B1(n29), .B2(n323), .A(n24), .ZN(n22) );
  NAND2_X1 U413 ( .A1(n96), .A2(n101), .ZN(n36) );
  OAI22_X1 U414 ( .A1(n328), .A2(n175), .B1(n174), .B2(n330), .ZN(n142) );
  OAI22_X1 U415 ( .A1(n328), .A2(n176), .B1(n175), .B2(n330), .ZN(n143) );
  OAI22_X1 U416 ( .A1(n329), .A2(n177), .B1(n176), .B2(n304), .ZN(n144) );
  OAI22_X1 U417 ( .A1(n328), .A2(n179), .B1(n178), .B2(n330), .ZN(n146) );
  INV_X1 U418 ( .A(n304), .ZN(n126) );
  XNOR2_X1 U419 ( .A(n278), .B(b[7]), .ZN(n182) );
  OAI22_X1 U420 ( .A1(n329), .A2(n178), .B1(n177), .B2(n304), .ZN(n145) );
  XNOR2_X1 U421 ( .A(n278), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U422 ( .A(n278), .B(b[6]), .ZN(n183) );
  OAI22_X1 U423 ( .A1(n221), .A2(n229), .B1(n181), .B2(n330), .ZN(n137) );
  OAI22_X1 U424 ( .A1(n221), .A2(n180), .B1(n179), .B2(n304), .ZN(n147) );
  XNOR2_X1 U425 ( .A(n278), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U426 ( .A(n278), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U427 ( .A(n334), .B(n278), .ZN(n189) );
  INV_X1 U428 ( .A(n234), .ZN(n230) );
  XOR2_X1 U429 ( .A(n234), .B(a[4]), .Z(n218) );
  XNOR2_X1 U430 ( .A(n282), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U431 ( .A(n278), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U432 ( .A(n233), .B(b[3]), .ZN(n177) );
  INV_X1 U433 ( .A(n317), .ZN(n73) );
  NAND2_X1 U434 ( .A1(n92), .A2(n95), .ZN(n31) );
  INV_X1 U435 ( .A(n320), .ZN(n75) );
  NOR2_X1 U436 ( .A1(n320), .A2(n44), .ZN(n39) );
  OAI21_X1 U437 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  NAND2_X1 U438 ( .A1(n102), .A2(n107), .ZN(n42) );
  INV_X1 U439 ( .A(n274), .ZN(n46) );
  OAI21_X1 U440 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  XOR2_X1 U441 ( .A(n7), .B(n318), .Z(product[6]) );
  AOI21_X1 U442 ( .B1(n326), .B2(n55), .A(n52), .ZN(n50) );
  XNOR2_X1 U443 ( .A(n234), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U444 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U445 ( .A(n276), .B(b[1]), .ZN(n197) );
  OAI22_X1 U446 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  NAND2_X1 U447 ( .A1(n171), .A2(n164), .ZN(n66) );
  INV_X1 U448 ( .A(n15), .ZN(n70) );
  OAI22_X1 U449 ( .A1(n182), .A2(n332), .B1(n182), .B2(n319), .ZN(n128) );
  OAI22_X1 U450 ( .A1(n332), .A2(n188), .B1(n187), .B2(n319), .ZN(n154) );
  OAI22_X1 U451 ( .A1(n332), .A2(n183), .B1(n182), .B2(n319), .ZN(n89) );
  OAI22_X1 U452 ( .A1(n332), .A2(n187), .B1(n186), .B2(n319), .ZN(n153) );
  OAI22_X1 U453 ( .A1(n333), .A2(n185), .B1(n184), .B2(n319), .ZN(n151) );
  OAI22_X1 U454 ( .A1(n332), .A2(n186), .B1(n185), .B2(n319), .ZN(n152) );
  OAI22_X1 U455 ( .A1(n333), .A2(n184), .B1(n183), .B2(n319), .ZN(n150) );
  INV_X1 U456 ( .A(n319), .ZN(n129) );
  OAI22_X1 U457 ( .A1(n222), .A2(n230), .B1(n190), .B2(n319), .ZN(n138) );
  OAI22_X1 U458 ( .A1(n222), .A2(n189), .B1(n188), .B2(n319), .ZN(n155) );
  OAI21_X1 U459 ( .B1(n315), .B2(n21), .A(n22), .ZN(n20) );
  XNOR2_X1 U460 ( .A(n307), .B(n1), .ZN(product[12]) );
  INV_X1 U461 ( .A(n301), .ZN(n37) );
  AOI21_X1 U462 ( .B1(n20), .B2(n325), .A(n17), .ZN(n15) );
  OAI22_X1 U463 ( .A1(n331), .A2(n193), .B1(n192), .B2(n327), .ZN(n158) );
  OAI22_X1 U464 ( .A1(n331), .A2(n195), .B1(n194), .B2(n327), .ZN(n160) );
  OAI22_X1 U465 ( .A1(n331), .A2(n194), .B1(n193), .B2(n327), .ZN(n159) );
  OAI22_X1 U466 ( .A1(n331), .A2(n196), .B1(n195), .B2(n327), .ZN(n161) );
  OAI22_X1 U467 ( .A1(n331), .A2(n231), .B1(n199), .B2(n327), .ZN(n139) );
  OAI22_X1 U468 ( .A1(n331), .A2(n197), .B1(n196), .B2(n327), .ZN(n162) );
  OAI22_X1 U469 ( .A1(n223), .A2(n192), .B1(n327), .B2(n191), .ZN(n99) );
  OAI22_X1 U470 ( .A1(n191), .A2(n223), .B1(n191), .B2(n327), .ZN(n131) );
  XNOR2_X1 U471 ( .A(n289), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U472 ( .A(n288), .B(b[6]), .ZN(n201) );
  INV_X1 U473 ( .A(n327), .ZN(n132) );
  OAI22_X1 U474 ( .A1(n331), .A2(n198), .B1(n197), .B2(n327), .ZN(n163) );
  XNOR2_X1 U475 ( .A(n288), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U476 ( .A(n289), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U477 ( .A(n334), .B(n289), .ZN(n207) );
  XNOR2_X1 U478 ( .A(n288), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U479 ( .A(n288), .B(b[3]), .ZN(n204) );
  INV_X1 U480 ( .A(n289), .ZN(n232) );
  XNOR2_X1 U481 ( .A(n288), .B(b[1]), .ZN(n206) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70,
         n73, n74, n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n128, n129, n131, n132, n134, n135, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n216, n217, n220, n221, n222, n223, n224, n225,
         n230, n231, n233, n234, n235, n236, n244, n274, n275, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n150), .B(n282), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n145), .B(n151), .CI(n100), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n166), .B(n159), .CI(n153), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n137), .B(n147), .CO(n111), .S(n112) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  OR2_X1 U237 ( .A1(n172), .A2(n140), .ZN(n274) );
  CLKBUF_X1 U238 ( .A(n31), .Z(n275) );
  AND3_X1 U239 ( .A1(n331), .A2(n330), .A3(n329), .ZN(product[15]) );
  CLKBUF_X1 U240 ( .A(n235), .Z(n277) );
  BUF_X1 U241 ( .A(n223), .Z(n287) );
  BUF_X1 U242 ( .A(n167), .Z(n278) );
  CLKBUF_X1 U243 ( .A(n45), .Z(n279) );
  OR2_X1 U244 ( .A1(n300), .A2(n301), .ZN(n222) );
  AOI21_X1 U245 ( .B1(n223), .B2(n343), .A(n191), .ZN(n131) );
  BUF_X1 U246 ( .A(n234), .Z(n280) );
  NAND2_X1 U247 ( .A1(n335), .A2(n336), .ZN(n281) );
  OAI22_X1 U248 ( .A1(n333), .A2(n192), .B1(n191), .B2(n343), .ZN(n282) );
  INV_X1 U249 ( .A(n233), .ZN(n283) );
  INV_X2 U250 ( .A(n283), .ZN(n284) );
  INV_X1 U251 ( .A(n126), .ZN(n285) );
  XNOR2_X1 U252 ( .A(n234), .B(a[6]), .ZN(n320) );
  OR2_X2 U253 ( .A1(n300), .A2(n301), .ZN(n286) );
  CLKBUF_X1 U254 ( .A(n236), .Z(n288) );
  CLKBUF_X1 U255 ( .A(n36), .Z(n289) );
  XOR2_X1 U256 ( .A(n167), .B(n148), .Z(n290) );
  XOR2_X1 U257 ( .A(n290), .B(n160), .Z(n116) );
  XOR2_X1 U258 ( .A(n119), .B(n154), .Z(n291) );
  XOR2_X1 U259 ( .A(n291), .B(n116), .Z(n114) );
  NAND2_X1 U260 ( .A1(n278), .A2(n148), .ZN(n292) );
  NAND2_X1 U261 ( .A1(n278), .A2(n160), .ZN(n293) );
  NAND2_X1 U262 ( .A1(n148), .A2(n160), .ZN(n294) );
  NAND3_X1 U263 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n115) );
  NAND2_X1 U264 ( .A1(n119), .A2(n154), .ZN(n295) );
  NAND2_X1 U265 ( .A1(n119), .A2(n116), .ZN(n296) );
  NAND2_X1 U266 ( .A1(n154), .A2(n116), .ZN(n297) );
  NAND3_X1 U267 ( .A1(n295), .A2(n296), .A3(n297), .ZN(n113) );
  NAND2_X1 U268 ( .A1(n220), .A2(n244), .ZN(n298) );
  NAND2_X1 U269 ( .A1(n220), .A2(n244), .ZN(n299) );
  NAND2_X1 U270 ( .A1(n220), .A2(n244), .ZN(n224) );
  XOR2_X1 U271 ( .A(n235), .B(a[4]), .Z(n300) );
  XNOR2_X1 U272 ( .A(n234), .B(a[4]), .ZN(n301) );
  INV_X1 U273 ( .A(n76), .ZN(n302) );
  XNOR2_X2 U274 ( .A(n236), .B(a[2]), .ZN(n343) );
  AOI21_X1 U275 ( .B1(n341), .B2(n55), .A(n52), .ZN(n303) );
  NOR2_X1 U276 ( .A1(n92), .A2(n95), .ZN(n304) );
  NOR2_X1 U277 ( .A1(n92), .A2(n95), .ZN(n30) );
  CLKBUF_X1 U278 ( .A(n221), .Z(n305) );
  NAND2_X1 U279 ( .A1(n217), .A2(n225), .ZN(n221) );
  CLKBUF_X1 U280 ( .A(n70), .Z(n306) );
  CLKBUF_X1 U281 ( .A(n40), .Z(n307) );
  NAND2_X1 U282 ( .A1(n236), .A2(n309), .ZN(n310) );
  NAND2_X1 U283 ( .A1(n308), .A2(n135), .ZN(n311) );
  NAND2_X1 U284 ( .A1(n310), .A2(n311), .ZN(n220) );
  INV_X1 U285 ( .A(n236), .ZN(n308) );
  INV_X1 U286 ( .A(n135), .ZN(n309) );
  NAND2_X1 U287 ( .A1(n235), .A2(n313), .ZN(n314) );
  NAND2_X1 U288 ( .A1(n312), .A2(a[2]), .ZN(n315) );
  NAND2_X1 U289 ( .A1(n314), .A2(n315), .ZN(n319) );
  INV_X1 U290 ( .A(n235), .ZN(n312) );
  INV_X1 U291 ( .A(a[2]), .ZN(n313) );
  INV_X1 U292 ( .A(n312), .ZN(n316) );
  XNOR2_X1 U293 ( .A(n317), .B(n323), .ZN(product[14]) );
  XNOR2_X1 U294 ( .A(n141), .B(n83), .ZN(n317) );
  CLKBUF_X1 U295 ( .A(n28), .Z(n318) );
  BUF_X2 U296 ( .A(n216), .Z(n352) );
  CLKBUF_X1 U297 ( .A(n234), .Z(n321) );
  NAND3_X1 U298 ( .A1(n327), .A2(n328), .A3(n326), .ZN(n322) );
  NAND3_X1 U299 ( .A1(n327), .A2(n328), .A3(n326), .ZN(n323) );
  CLKBUF_X1 U300 ( .A(n20), .Z(n324) );
  XOR2_X1 U301 ( .A(n85), .B(n84), .Z(n325) );
  XOR2_X1 U302 ( .A(n325), .B(n306), .Z(product[13]) );
  NAND2_X1 U303 ( .A1(n85), .A2(n84), .ZN(n326) );
  NAND2_X1 U304 ( .A1(n70), .A2(n85), .ZN(n327) );
  NAND2_X1 U305 ( .A1(n70), .A2(n84), .ZN(n328) );
  NAND3_X1 U306 ( .A1(n328), .A2(n327), .A3(n326), .ZN(n14) );
  NAND2_X1 U307 ( .A1(n141), .A2(n83), .ZN(n329) );
  NAND2_X1 U308 ( .A1(n141), .A2(n14), .ZN(n330) );
  NAND2_X1 U309 ( .A1(n83), .A2(n322), .ZN(n331) );
  NOR2_X2 U310 ( .A1(n114), .A2(n117), .ZN(n48) );
  CLKBUF_X1 U311 ( .A(n29), .Z(n332) );
  AOI21_X1 U312 ( .B1(n341), .B2(n55), .A(n52), .ZN(n50) );
  NAND2_X1 U313 ( .A1(n336), .A2(n335), .ZN(n333) );
  AOI21_X1 U314 ( .B1(n39), .B2(n348), .A(n307), .ZN(n334) );
  NAND2_X1 U315 ( .A1(n336), .A2(n319), .ZN(n223) );
  NOR2_X1 U316 ( .A1(n108), .A2(n113), .ZN(n44) );
  NAND2_X1 U317 ( .A1(n108), .A2(n113), .ZN(n45) );
  OR2_X1 U318 ( .A1(n88), .A2(n91), .ZN(n338) );
  XOR2_X1 U319 ( .A(n235), .B(a[2]), .Z(n335) );
  XNOR2_X1 U320 ( .A(n236), .B(a[2]), .ZN(n336) );
  XNOR2_X1 U321 ( .A(n37), .B(n4), .ZN(product[9]) );
  INV_X1 U322 ( .A(n35), .ZN(n74) );
  INV_X1 U323 ( .A(n66), .ZN(n64) );
  INV_X1 U324 ( .A(n26), .ZN(n24) );
  OAI21_X1 U325 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  NAND2_X1 U326 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U327 ( .A(n48), .ZN(n77) );
  NAND2_X1 U328 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U329 ( .A(n60), .ZN(n80) );
  NAND2_X1 U330 ( .A1(n340), .A2(n19), .ZN(n1) );
  XOR2_X1 U331 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U332 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U333 ( .A(n56), .ZN(n79) );
  XOR2_X1 U334 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U335 ( .A1(n73), .A2(n275), .ZN(n3) );
  AOI21_X1 U336 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U337 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U338 ( .A1(n76), .A2(n279), .ZN(n6) );
  INV_X1 U339 ( .A(n44), .ZN(n76) );
  XOR2_X1 U340 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U341 ( .A1(n338), .A2(n26), .ZN(n2) );
  XNOR2_X1 U342 ( .A(n8), .B(n55), .ZN(product[5]) );
  XNOR2_X1 U343 ( .A(n43), .B(n5), .ZN(product[8]) );
  OAI21_X1 U344 ( .B1(n46), .B2(n302), .A(n279), .ZN(n43) );
  XNOR2_X1 U345 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U346 ( .A1(n339), .A2(n66), .ZN(n11) );
  INV_X1 U347 ( .A(n59), .ZN(n58) );
  INV_X1 U348 ( .A(n19), .ZN(n17) );
  XNOR2_X1 U349 ( .A(n104), .B(n337), .ZN(n102) );
  XNOR2_X1 U350 ( .A(n106), .B(n109), .ZN(n337) );
  NOR2_X1 U351 ( .A1(n122), .A2(n123), .ZN(n56) );
  OR2_X1 U352 ( .A1(n158), .A2(n146), .ZN(n105) );
  NAND2_X1 U353 ( .A1(n124), .A2(n139), .ZN(n61) );
  INV_X1 U354 ( .A(n83), .ZN(n84) );
  NAND2_X1 U355 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U356 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U357 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U358 ( .A1(n122), .A2(n123), .ZN(n57) );
  INV_X1 U359 ( .A(n69), .ZN(n67) );
  OR2_X1 U360 ( .A1(n171), .A2(n164), .ZN(n339) );
  OR2_X1 U361 ( .A1(n87), .A2(n86), .ZN(n340) );
  OR2_X1 U362 ( .A1(n118), .A2(n121), .ZN(n341) );
  OR2_X1 U363 ( .A1(n352), .A2(n231), .ZN(n199) );
  AND2_X1 U364 ( .A1(n352), .A2(n126), .ZN(n148) );
  INV_X1 U365 ( .A(n128), .ZN(n149) );
  INV_X1 U366 ( .A(n89), .ZN(n90) );
  AND2_X1 U367 ( .A1(n352), .A2(n129), .ZN(n156) );
  OAI22_X1 U368 ( .A1(n299), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OR2_X1 U369 ( .A1(n352), .A2(n230), .ZN(n190) );
  OAI22_X1 U370 ( .A1(n298), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  INV_X1 U371 ( .A(n134), .ZN(n165) );
  OAI22_X1 U372 ( .A1(n200), .A2(n298), .B1(n200), .B2(n244), .ZN(n134) );
  INV_X1 U373 ( .A(n125), .ZN(n141) );
  OR2_X1 U374 ( .A1(n352), .A2(n283), .ZN(n181) );
  AND2_X1 U375 ( .A1(n274), .A2(n69), .ZN(product[1]) );
  AND2_X1 U376 ( .A1(n352), .A2(n132), .ZN(n164) );
  OR2_X1 U377 ( .A1(n352), .A2(n308), .ZN(n208) );
  OAI22_X1 U378 ( .A1(n299), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  AND2_X1 U379 ( .A1(n352), .A2(n135), .ZN(product[0]) );
  NOR2_X1 U380 ( .A1(n124), .A2(n139), .ZN(n60) );
  NAND2_X1 U381 ( .A1(n341), .A2(n54), .ZN(n8) );
  INV_X1 U382 ( .A(n54), .ZN(n52) );
  XNOR2_X1 U383 ( .A(n234), .B(a[6]), .ZN(n225) );
  XNOR2_X1 U384 ( .A(n284), .B(b[7]), .ZN(n173) );
  XNOR2_X1 U385 ( .A(n284), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U386 ( .A(n284), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U387 ( .A(n284), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U388 ( .A(n284), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U389 ( .A(n284), .B(b[2]), .ZN(n178) );
  XOR2_X1 U390 ( .A(n233), .B(a[6]), .Z(n217) );
  XNOR2_X2 U391 ( .A(n235), .B(a[4]), .ZN(n347) );
  OAI22_X1 U392 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U393 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI21_X1 U394 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  INV_X1 U395 ( .A(n289), .ZN(n34) );
  NAND2_X1 U396 ( .A1(n74), .A2(n289), .ZN(n4) );
  INV_X1 U397 ( .A(n99), .ZN(n100) );
  INV_X1 U398 ( .A(n131), .ZN(n157) );
  NAND2_X1 U399 ( .A1(n104), .A2(n106), .ZN(n344) );
  NAND2_X1 U400 ( .A1(n104), .A2(n109), .ZN(n345) );
  NAND2_X1 U401 ( .A1(n106), .A2(n109), .ZN(n346) );
  NAND3_X1 U402 ( .A1(n344), .A2(n345), .A3(n346), .ZN(n101) );
  XNOR2_X1 U403 ( .A(n158), .B(n146), .ZN(n106) );
  XOR2_X1 U404 ( .A(n10), .B(n62), .Z(product[3]) );
  OAI21_X1 U405 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  AOI21_X1 U406 ( .B1(n339), .B2(n67), .A(n64), .ZN(n62) );
  NAND2_X1 U407 ( .A1(n172), .A2(n140), .ZN(n69) );
  NAND2_X1 U408 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U409 ( .B1(n48), .B2(n303), .A(n49), .ZN(n348) );
  NOR2_X1 U410 ( .A1(n107), .A2(n102), .ZN(n349) );
  OR2_X1 U411 ( .A1(n221), .A2(n180), .ZN(n350) );
  OR2_X1 U412 ( .A1(n179), .A2(n320), .ZN(n351) );
  NAND2_X1 U413 ( .A1(n350), .A2(n351), .ZN(n147) );
  NOR2_X1 U414 ( .A1(n102), .A2(n107), .ZN(n41) );
  XNOR2_X1 U415 ( .A(n216), .B(n233), .ZN(n180) );
  NAND2_X1 U416 ( .A1(n96), .A2(n101), .ZN(n36) );
  NOR2_X1 U417 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U418 ( .A1(n118), .A2(n121), .ZN(n54) );
  AOI21_X1 U419 ( .B1(n37), .B2(n318), .A(n332), .ZN(n27) );
  NAND2_X1 U420 ( .A1(n28), .A2(n338), .ZN(n21) );
  NOR2_X1 U421 ( .A1(n35), .A2(n304), .ZN(n28) );
  OAI22_X1 U422 ( .A1(n298), .A2(n308), .B1(n208), .B2(n244), .ZN(n140) );
  AOI21_X1 U423 ( .B1(n29), .B2(n338), .A(n24), .ZN(n22) );
  OAI22_X1 U424 ( .A1(n299), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  NAND2_X1 U425 ( .A1(n171), .A2(n164), .ZN(n66) );
  XNOR2_X1 U426 ( .A(n236), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U427 ( .A(n236), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U428 ( .A(n288), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U429 ( .A(n352), .B(n288), .ZN(n207) );
  XNOR2_X1 U430 ( .A(n236), .B(b[3]), .ZN(n204) );
  XNOR2_X1 U431 ( .A(n236), .B(b[7]), .ZN(n200) );
  OAI21_X1 U432 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  OAI22_X1 U433 ( .A1(n182), .A2(n286), .B1(n182), .B2(n347), .ZN(n128) );
  OAI22_X1 U434 ( .A1(n286), .A2(n188), .B1(n187), .B2(n347), .ZN(n154) );
  OAI22_X1 U435 ( .A1(n286), .A2(n183), .B1(n182), .B2(n347), .ZN(n89) );
  OAI22_X1 U436 ( .A1(n222), .A2(n184), .B1(n183), .B2(n347), .ZN(n150) );
  OAI22_X1 U437 ( .A1(n286), .A2(n187), .B1(n186), .B2(n347), .ZN(n153) );
  OAI22_X1 U438 ( .A1(n286), .A2(n186), .B1(n185), .B2(n347), .ZN(n152) );
  INV_X1 U439 ( .A(n347), .ZN(n129) );
  OAI22_X1 U440 ( .A1(n286), .A2(n185), .B1(n184), .B2(n347), .ZN(n151) );
  XNOR2_X1 U441 ( .A(n277), .B(b[3]), .ZN(n195) );
  OAI22_X1 U442 ( .A1(n222), .A2(n230), .B1(n190), .B2(n347), .ZN(n138) );
  OAI22_X1 U443 ( .A1(n222), .A2(n189), .B1(n188), .B2(n347), .ZN(n155) );
  XNOR2_X1 U444 ( .A(n277), .B(b[4]), .ZN(n194) );
  INV_X1 U445 ( .A(n316), .ZN(n231) );
  XNOR2_X1 U446 ( .A(n235), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U447 ( .A(n316), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U448 ( .A(n352), .B(n316), .ZN(n198) );
  XNOR2_X1 U449 ( .A(n235), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U450 ( .A(b[7]), .B(n235), .ZN(n191) );
  INV_X1 U451 ( .A(n304), .ZN(n73) );
  NAND2_X1 U452 ( .A1(n92), .A2(n95), .ZN(n31) );
  INV_X1 U453 ( .A(n348), .ZN(n46) );
  AOI21_X1 U454 ( .B1(n39), .B2(n47), .A(n40), .ZN(n38) );
  OAI21_X1 U455 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  XOR2_X1 U456 ( .A(n7), .B(n303), .Z(product[6]) );
  INV_X1 U457 ( .A(n349), .ZN(n75) );
  OAI22_X1 U458 ( .A1(n173), .A2(n305), .B1(n173), .B2(n285), .ZN(n125) );
  OAI22_X1 U459 ( .A1(n305), .A2(n174), .B1(n173), .B2(n285), .ZN(n83) );
  NOR2_X1 U460 ( .A1(n349), .A2(n44), .ZN(n39) );
  OAI21_X1 U461 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  NAND2_X1 U462 ( .A1(n102), .A2(n107), .ZN(n42) );
  OAI22_X1 U463 ( .A1(n305), .A2(n175), .B1(n174), .B2(n285), .ZN(n142) );
  OAI22_X1 U464 ( .A1(n305), .A2(n176), .B1(n175), .B2(n285), .ZN(n143) );
  OAI22_X1 U465 ( .A1(n305), .A2(n177), .B1(n176), .B2(n285), .ZN(n144) );
  XNOR2_X1 U466 ( .A(n321), .B(b[7]), .ZN(n182) );
  OAI22_X1 U467 ( .A1(n221), .A2(n178), .B1(n177), .B2(n320), .ZN(n145) );
  INV_X1 U468 ( .A(n320), .ZN(n126) );
  OAI22_X1 U469 ( .A1(n221), .A2(n179), .B1(n178), .B2(n285), .ZN(n146) );
  XNOR2_X1 U470 ( .A(n280), .B(b[5]), .ZN(n184) );
  OAI22_X1 U471 ( .A1(n221), .A2(n283), .B1(n181), .B2(n320), .ZN(n137) );
  XNOR2_X1 U472 ( .A(n280), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U473 ( .A(n280), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U474 ( .A(n280), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U475 ( .A(n321), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U476 ( .A(n352), .B(n321), .ZN(n189) );
  INV_X1 U477 ( .A(n234), .ZN(n230) );
  XNOR2_X1 U478 ( .A(n288), .B(b[2]), .ZN(n205) );
  INV_X1 U479 ( .A(n15), .ZN(n70) );
  OAI22_X1 U480 ( .A1(n298), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  XNOR2_X1 U481 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U482 ( .A(n280), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U483 ( .A(b[1]), .B(n277), .ZN(n197) );
  XNOR2_X1 U484 ( .A(n236), .B(b[1]), .ZN(n206) );
  XNOR2_X1 U485 ( .A(n324), .B(n1), .ZN(product[12]) );
  INV_X1 U486 ( .A(n334), .ZN(n37) );
  AOI21_X1 U487 ( .B1(n20), .B2(n340), .A(n17), .ZN(n15) );
  OAI22_X1 U488 ( .A1(n281), .A2(n193), .B1(n192), .B2(n343), .ZN(n158) );
  OAI22_X1 U489 ( .A1(n223), .A2(n195), .B1(n194), .B2(n343), .ZN(n160) );
  OAI22_X1 U490 ( .A1(n194), .A2(n333), .B1(n193), .B2(n343), .ZN(n159) );
  OAI22_X1 U491 ( .A1(n287), .A2(n196), .B1(n195), .B2(n343), .ZN(n161) );
  OAI22_X1 U492 ( .A1(n287), .A2(n231), .B1(n199), .B2(n343), .ZN(n139) );
  OAI22_X1 U493 ( .A1(n287), .A2(n197), .B1(n196), .B2(n343), .ZN(n162) );
  OAI22_X1 U494 ( .A1(n281), .A2(n192), .B1(n191), .B2(n343), .ZN(n99) );
  INV_X1 U495 ( .A(n343), .ZN(n132) );
  OAI22_X1 U496 ( .A1(n281), .A2(n198), .B1(n197), .B2(n343), .ZN(n163) );
  INV_X2 U497 ( .A(n135), .ZN(n244) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70,
         n74, n75, n76, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n129, n132, n134, n135, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n216,
         n217, n218, n219, n221, n222, n223, n224, n225, n226, n227, n229,
         n230, n231, n232, n233, n234, n235, n236, n244, n274, n275, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U103 ( .A(n145), .B(n151), .CI(n100), .CO(n97), .S(n98) );
  FA_X1 U105 ( .A(n109), .B(n106), .CI(n104), .CO(n101), .S(n102) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n166), .B(n153), .CI(n159), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  BUF_X1 U237 ( .A(n234), .Z(n304) );
  BUF_X1 U238 ( .A(n234), .Z(n330) );
  BUF_X2 U239 ( .A(n235), .Z(n342) );
  BUF_X2 U240 ( .A(n216), .Z(n292) );
  AND2_X1 U241 ( .A1(n327), .A2(n328), .ZN(n274) );
  OR2_X1 U242 ( .A1(n92), .A2(n95), .ZN(n275) );
  AND2_X1 U243 ( .A1(n337), .A2(n69), .ZN(product[1]) );
  CLKBUF_X3 U244 ( .A(n225), .Z(n335) );
  XNOR2_X1 U245 ( .A(n290), .B(b[7]), .ZN(n277) );
  CLKBUF_X1 U246 ( .A(n45), .Z(n278) );
  XOR2_X1 U247 ( .A(n103), .B(n105), .Z(n279) );
  XOR2_X1 U248 ( .A(n98), .B(n279), .Z(n96) );
  NAND2_X1 U249 ( .A1(n98), .A2(n103), .ZN(n280) );
  NAND2_X1 U250 ( .A1(n98), .A2(n105), .ZN(n281) );
  NAND2_X1 U251 ( .A1(n103), .A2(n105), .ZN(n282) );
  NAND3_X1 U252 ( .A1(n280), .A2(n281), .A3(n282), .ZN(n95) );
  OR2_X1 U253 ( .A1(n114), .A2(n117), .ZN(n283) );
  NOR2_X1 U254 ( .A1(n92), .A2(n95), .ZN(n284) );
  CLKBUF_X1 U255 ( .A(n28), .Z(n285) );
  NOR2_X1 U256 ( .A1(n92), .A2(n95), .ZN(n30) );
  CLKBUF_X1 U257 ( .A(n55), .Z(n286) );
  CLKBUF_X1 U258 ( .A(n217), .Z(n287) );
  BUF_X2 U259 ( .A(n226), .Z(n349) );
  BUF_X2 U260 ( .A(n226), .Z(n348) );
  NAND2_X1 U261 ( .A1(n219), .A2(n227), .ZN(n288) );
  NAND2_X1 U262 ( .A1(n219), .A2(n227), .ZN(n289) );
  NAND2_X1 U263 ( .A1(n219), .A2(n227), .ZN(n223) );
  BUF_X2 U264 ( .A(n236), .Z(n290) );
  INV_X1 U265 ( .A(n76), .ZN(n291) );
  XNOR2_X1 U266 ( .A(n341), .B(a[4]), .ZN(n293) );
  BUF_X1 U267 ( .A(n235), .Z(n341) );
  CLKBUF_X1 U268 ( .A(n47), .Z(n294) );
  CLKBUF_X1 U269 ( .A(n288), .Z(n295) );
  INV_X1 U270 ( .A(n229), .ZN(n296) );
  CLKBUF_X1 U271 ( .A(n50), .Z(n297) );
  AOI21_X1 U272 ( .B1(n336), .B2(n55), .A(n52), .ZN(n50) );
  CLKBUF_X1 U273 ( .A(n227), .Z(n344) );
  NAND2_X1 U274 ( .A1(n342), .A2(n299), .ZN(n300) );
  NAND2_X1 U275 ( .A1(n298), .A2(a[2]), .ZN(n301) );
  NAND2_X1 U276 ( .A1(n301), .A2(n300), .ZN(n219) );
  INV_X1 U277 ( .A(n342), .ZN(n298) );
  INV_X1 U278 ( .A(a[2]), .ZN(n299) );
  XNOR2_X1 U279 ( .A(n234), .B(a[6]), .ZN(n302) );
  XNOR2_X1 U280 ( .A(n234), .B(a[6]), .ZN(n225) );
  CLKBUF_X1 U281 ( .A(n221), .Z(n303) );
  NAND3_X1 U282 ( .A1(n313), .A2(n312), .A3(n311), .ZN(n305) );
  XNOR2_X1 U283 ( .A(n305), .B(n306), .ZN(product[14]) );
  XNOR2_X1 U284 ( .A(n141), .B(n83), .ZN(n306) );
  AND3_X1 U285 ( .A1(n315), .A2(n316), .A3(n314), .ZN(product[15]) );
  CLKBUF_X1 U286 ( .A(n70), .Z(n308) );
  XNOR2_X1 U287 ( .A(n309), .B(n274), .ZN(n94) );
  XNOR2_X1 U288 ( .A(n150), .B(n333), .ZN(n309) );
  XOR2_X1 U289 ( .A(n85), .B(n84), .Z(n310) );
  XOR2_X1 U290 ( .A(n310), .B(n308), .Z(product[13]) );
  NAND2_X1 U291 ( .A1(n85), .A2(n84), .ZN(n311) );
  NAND2_X1 U292 ( .A1(n70), .A2(n85), .ZN(n312) );
  NAND2_X1 U293 ( .A1(n70), .A2(n84), .ZN(n313) );
  NAND3_X1 U294 ( .A1(n312), .A2(n313), .A3(n311), .ZN(n14) );
  NAND2_X1 U295 ( .A1(n141), .A2(n83), .ZN(n314) );
  NAND2_X1 U296 ( .A1(n305), .A2(n141), .ZN(n315) );
  NAND2_X1 U297 ( .A1(n83), .A2(n14), .ZN(n316) );
  CLKBUF_X1 U298 ( .A(n39), .Z(n317) );
  CLKBUF_X1 U299 ( .A(n346), .Z(n318) );
  XNOR2_X1 U300 ( .A(n319), .B(n94), .ZN(n92) );
  XNOR2_X1 U301 ( .A(n97), .B(n144), .ZN(n319) );
  CLKBUF_X1 U302 ( .A(n40), .Z(n320) );
  NAND2_X1 U303 ( .A1(n150), .A2(n333), .ZN(n321) );
  NAND2_X1 U304 ( .A1(n150), .A2(n274), .ZN(n322) );
  NAND2_X1 U305 ( .A1(n274), .A2(n333), .ZN(n323) );
  NAND3_X1 U306 ( .A1(n321), .A2(n322), .A3(n323), .ZN(n93) );
  NAND2_X1 U307 ( .A1(n97), .A2(n144), .ZN(n324) );
  NAND2_X1 U308 ( .A1(n97), .A2(n94), .ZN(n325) );
  NAND2_X1 U309 ( .A1(n144), .A2(n94), .ZN(n326) );
  NAND3_X1 U310 ( .A1(n324), .A2(n325), .A3(n326), .ZN(n91) );
  OR2_X1 U311 ( .A1(n288), .A2(n191), .ZN(n327) );
  OR2_X1 U312 ( .A1(n191), .A2(n344), .ZN(n328) );
  OR2_X2 U313 ( .A1(n329), .A2(n135), .ZN(n224) );
  XNOR2_X1 U314 ( .A(n236), .B(n135), .ZN(n329) );
  INV_X1 U315 ( .A(n135), .ZN(n244) );
  CLKBUF_X1 U316 ( .A(n42), .Z(n331) );
  CLKBUF_X1 U317 ( .A(n20), .Z(n332) );
  OAI22_X1 U318 ( .A1(n288), .A2(n192), .B1(n191), .B2(n344), .ZN(n333) );
  AOI21_X1 U319 ( .B1(n317), .B2(n294), .A(n320), .ZN(n334) );
  NOR2_X1 U320 ( .A1(n108), .A2(n113), .ZN(n44) );
  NAND2_X1 U321 ( .A1(n108), .A2(n113), .ZN(n45) );
  OR2_X1 U322 ( .A1(n118), .A2(n121), .ZN(n336) );
  OR2_X1 U323 ( .A1(n172), .A2(n140), .ZN(n337) );
  INV_X1 U324 ( .A(n35), .ZN(n74) );
  XNOR2_X1 U325 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U326 ( .A1(n74), .A2(n36), .ZN(n4) );
  INV_X1 U327 ( .A(n36), .ZN(n34) );
  INV_X1 U328 ( .A(n66), .ZN(n64) );
  INV_X1 U329 ( .A(n26), .ZN(n24) );
  OAI21_X1 U330 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  NOR2_X1 U331 ( .A1(n96), .A2(n101), .ZN(n35) );
  INV_X1 U332 ( .A(n54), .ZN(n52) );
  NAND2_X1 U333 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U334 ( .A(n60), .ZN(n80) );
  NAND2_X1 U335 ( .A1(n96), .A2(n101), .ZN(n36) );
  NAND2_X1 U336 ( .A1(n340), .A2(n19), .ZN(n1) );
  XOR2_X1 U337 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U338 ( .A1(n275), .A2(n31), .ZN(n3) );
  AOI21_X1 U339 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U340 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U341 ( .A1(n76), .A2(n278), .ZN(n6) );
  INV_X1 U342 ( .A(n44), .ZN(n76) );
  XOR2_X1 U343 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U344 ( .A1(n338), .A2(n26), .ZN(n2) );
  NOR2_X1 U345 ( .A1(n35), .A2(n30), .ZN(n28) );
  XNOR2_X1 U346 ( .A(n43), .B(n5), .ZN(product[8]) );
  OAI21_X1 U347 ( .B1(n46), .B2(n291), .A(n278), .ZN(n43) );
  XNOR2_X1 U348 ( .A(n8), .B(n286), .ZN(product[5]) );
  NAND2_X1 U349 ( .A1(n336), .A2(n54), .ZN(n8) );
  XNOR2_X1 U350 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U351 ( .A1(n339), .A2(n66), .ZN(n11) );
  INV_X1 U352 ( .A(n59), .ZN(n58) );
  NAND2_X1 U353 ( .A1(n283), .A2(n49), .ZN(n7) );
  XOR2_X1 U354 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U355 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U356 ( .A(n56), .ZN(n79) );
  INV_X1 U357 ( .A(n19), .ZN(n17) );
  OR2_X1 U358 ( .A1(n158), .A2(n146), .ZN(n105) );
  XNOR2_X1 U359 ( .A(n158), .B(n146), .ZN(n106) );
  NOR2_X1 U360 ( .A1(n122), .A2(n123), .ZN(n56) );
  NOR2_X1 U361 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U362 ( .A(n69), .ZN(n67) );
  INV_X1 U363 ( .A(n83), .ZN(n84) );
  OR2_X2 U364 ( .A1(n88), .A2(n91), .ZN(n338) );
  NAND2_X1 U365 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U366 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U367 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U368 ( .A1(n122), .A2(n123), .ZN(n57) );
  OR2_X1 U369 ( .A1(n171), .A2(n164), .ZN(n339) );
  NAND2_X1 U370 ( .A1(n92), .A2(n95), .ZN(n31) );
  OR2_X1 U371 ( .A1(n87), .A2(n86), .ZN(n340) );
  AND2_X1 U372 ( .A1(n292), .A2(n132), .ZN(n164) );
  INV_X1 U373 ( .A(n128), .ZN(n149) );
  OR2_X1 U374 ( .A1(n292), .A2(n231), .ZN(n199) );
  AND2_X1 U375 ( .A1(n292), .A2(n129), .ZN(n156) );
  INV_X1 U376 ( .A(n89), .ZN(n90) );
  INV_X1 U377 ( .A(n134), .ZN(n165) );
  AND2_X1 U378 ( .A1(n292), .A2(n126), .ZN(n148) );
  INV_X1 U379 ( .A(n125), .ZN(n141) );
  OR2_X1 U380 ( .A1(n216), .A2(n229), .ZN(n181) );
  OR2_X1 U381 ( .A1(n292), .A2(n230), .ZN(n190) );
  OR2_X1 U382 ( .A1(n292), .A2(n232), .ZN(n208) );
  XNOR2_X1 U383 ( .A(n296), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U384 ( .A(n296), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U385 ( .A(n296), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U386 ( .A(n296), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U387 ( .A(n216), .B(n233), .ZN(n180) );
  INV_X1 U388 ( .A(n233), .ZN(n229) );
  AND2_X1 U389 ( .A1(n292), .A2(n135), .ZN(product[0]) );
  NAND2_X1 U390 ( .A1(n124), .A2(n139), .ZN(n61) );
  NAND2_X1 U391 ( .A1(n75), .A2(n331), .ZN(n5) );
  OAI22_X1 U392 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  OAI22_X1 U393 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U394 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U395 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  OAI22_X1 U396 ( .A1(n224), .A2(n201), .B1(n277), .B2(n244), .ZN(n166) );
  OAI22_X1 U397 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  NAND2_X1 U398 ( .A1(n218), .A2(n293), .ZN(n343) );
  NAND2_X1 U399 ( .A1(n218), .A2(n293), .ZN(n222) );
  CLKBUF_X1 U400 ( .A(n227), .Z(n345) );
  XNOR2_X1 U401 ( .A(n236), .B(a[2]), .ZN(n227) );
  NOR2_X1 U402 ( .A1(n107), .A2(n102), .ZN(n346) );
  NAND2_X1 U403 ( .A1(n287), .A2(n335), .ZN(n347) );
  NOR2_X1 U404 ( .A1(n102), .A2(n107), .ZN(n41) );
  NAND2_X1 U405 ( .A1(n217), .A2(n225), .ZN(n221) );
  NAND2_X1 U406 ( .A1(n172), .A2(n140), .ZN(n69) );
  AOI21_X1 U407 ( .B1(n37), .B2(n285), .A(n29), .ZN(n27) );
  INV_X1 U408 ( .A(n99), .ZN(n100) );
  OAI22_X1 U409 ( .A1(n277), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  XNOR2_X1 U410 ( .A(n341), .B(a[4]), .ZN(n226) );
  XNOR2_X1 U411 ( .A(n296), .B(b[3]), .ZN(n177) );
  AOI21_X1 U412 ( .B1(n339), .B2(n67), .A(n64), .ZN(n62) );
  NOR2_X1 U413 ( .A1(n124), .A2(n139), .ZN(n60) );
  OAI22_X1 U414 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  XOR2_X1 U415 ( .A(n233), .B(a[6]), .Z(n217) );
  OAI22_X1 U416 ( .A1(n182), .A2(n343), .B1(n182), .B2(n348), .ZN(n128) );
  OAI22_X1 U417 ( .A1(n343), .A2(n188), .B1(n187), .B2(n349), .ZN(n154) );
  OAI22_X1 U418 ( .A1(n343), .A2(n183), .B1(n182), .B2(n348), .ZN(n89) );
  OAI22_X1 U419 ( .A1(n343), .A2(n185), .B1(n184), .B2(n348), .ZN(n151) );
  OAI22_X1 U420 ( .A1(n343), .A2(n184), .B1(n183), .B2(n349), .ZN(n150) );
  OAI22_X1 U421 ( .A1(n343), .A2(n186), .B1(n185), .B2(n349), .ZN(n152) );
  OAI22_X1 U422 ( .A1(n222), .A2(n187), .B1(n186), .B2(n349), .ZN(n153) );
  OAI22_X1 U423 ( .A1(n222), .A2(n230), .B1(n190), .B2(n348), .ZN(n138) );
  OAI22_X1 U424 ( .A1(n222), .A2(n189), .B1(n188), .B2(n349), .ZN(n155) );
  INV_X1 U425 ( .A(n348), .ZN(n129) );
  XOR2_X1 U426 ( .A(n10), .B(n62), .Z(product[3]) );
  OAI21_X1 U427 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  NAND2_X1 U428 ( .A1(n171), .A2(n164), .ZN(n66) );
  XNOR2_X1 U429 ( .A(n233), .B(b[1]), .ZN(n179) );
  INV_X1 U430 ( .A(n318), .ZN(n75) );
  NOR2_X1 U431 ( .A1(n346), .A2(n44), .ZN(n39) );
  OAI21_X1 U432 ( .B1(n284), .B2(n36), .A(n31), .ZN(n29) );
  NAND2_X1 U433 ( .A1(n118), .A2(n121), .ZN(n54) );
  XNOR2_X1 U434 ( .A(n296), .B(b[7]), .ZN(n173) );
  NAND2_X1 U435 ( .A1(n102), .A2(n107), .ZN(n42) );
  XNOR2_X1 U436 ( .A(n330), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U437 ( .A(n304), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U438 ( .A(n330), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U439 ( .A(n304), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U440 ( .A(n330), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U441 ( .A(n304), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U442 ( .A(n292), .B(n304), .ZN(n189) );
  INV_X1 U443 ( .A(n234), .ZN(n230) );
  XNOR2_X1 U444 ( .A(n330), .B(b[1]), .ZN(n188) );
  XOR2_X1 U445 ( .A(n234), .B(a[4]), .Z(n218) );
  NAND2_X1 U446 ( .A1(n28), .A2(n338), .ZN(n21) );
  OAI22_X1 U447 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI21_X1 U448 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U449 ( .B1(n29), .B2(n338), .A(n24), .ZN(n22) );
  OAI21_X1 U450 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  XOR2_X1 U451 ( .A(n7), .B(n297), .Z(product[6]) );
  INV_X1 U452 ( .A(n294), .ZN(n46) );
  AOI21_X1 U453 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U454 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  XNOR2_X1 U455 ( .A(n342), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U456 ( .A(n342), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U457 ( .A(n342), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U458 ( .A(n342), .B(b[2]), .ZN(n196) );
  INV_X1 U459 ( .A(n342), .ZN(n231) );
  XNOR2_X1 U460 ( .A(n342), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U461 ( .A(n342), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U462 ( .A(n292), .B(n342), .ZN(n198) );
  XNOR2_X1 U463 ( .A(n342), .B(b[1]), .ZN(n197) );
  INV_X1 U464 ( .A(n15), .ZN(n70) );
  OAI22_X1 U465 ( .A1(n173), .A2(n347), .B1(n173), .B2(n335), .ZN(n125) );
  OAI22_X1 U466 ( .A1(n347), .A2(n174), .B1(n173), .B2(n335), .ZN(n83) );
  OAI22_X1 U467 ( .A1(n347), .A2(n175), .B1(n174), .B2(n335), .ZN(n142) );
  OAI22_X1 U468 ( .A1(n347), .A2(n176), .B1(n175), .B2(n335), .ZN(n143) );
  OAI22_X1 U469 ( .A1(n347), .A2(n177), .B1(n176), .B2(n335), .ZN(n144) );
  OAI22_X1 U470 ( .A1(n347), .A2(n179), .B1(n178), .B2(n335), .ZN(n146) );
  OAI22_X1 U471 ( .A1(n303), .A2(n178), .B1(n177), .B2(n335), .ZN(n145) );
  INV_X1 U472 ( .A(n302), .ZN(n126) );
  OAI22_X1 U473 ( .A1(n221), .A2(n229), .B1(n181), .B2(n302), .ZN(n137) );
  OAI22_X1 U474 ( .A1(n221), .A2(n180), .B1(n179), .B2(n302), .ZN(n147) );
  XNOR2_X1 U475 ( .A(n332), .B(n1), .ZN(product[12]) );
  INV_X1 U476 ( .A(n334), .ZN(n37) );
  AOI21_X1 U477 ( .B1(n20), .B2(n340), .A(n17), .ZN(n15) );
  OAI22_X1 U478 ( .A1(n289), .A2(n193), .B1(n192), .B2(n344), .ZN(n158) );
  OAI22_X1 U479 ( .A1(n289), .A2(n195), .B1(n194), .B2(n344), .ZN(n160) );
  OAI22_X1 U480 ( .A1(n223), .A2(n194), .B1(n193), .B2(n345), .ZN(n159) );
  OAI22_X1 U481 ( .A1(n288), .A2(n196), .B1(n195), .B2(n344), .ZN(n161) );
  OAI22_X1 U482 ( .A1(n295), .A2(n231), .B1(n199), .B2(n344), .ZN(n139) );
  OAI22_X1 U483 ( .A1(n289), .A2(n197), .B1(n196), .B2(n345), .ZN(n162) );
  OAI22_X1 U484 ( .A1(n223), .A2(n192), .B1(n191), .B2(n344), .ZN(n99) );
  XNOR2_X1 U485 ( .A(n290), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U486 ( .A(n290), .B(b[6]), .ZN(n201) );
  INV_X1 U487 ( .A(n345), .ZN(n132) );
  OAI22_X1 U488 ( .A1(n288), .A2(n198), .B1(n197), .B2(n345), .ZN(n163) );
  XNOR2_X1 U489 ( .A(n290), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U490 ( .A(n290), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U491 ( .A(n292), .B(n290), .ZN(n207) );
  XNOR2_X1 U492 ( .A(n290), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U493 ( .A(n290), .B(b[3]), .ZN(n204) );
  INV_X1 U494 ( .A(n290), .ZN(n232) );
  XNOR2_X1 U495 ( .A(n290), .B(b[1]), .ZN(n206) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70,
         n74, n75, n76, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n129, n131, n134, n135, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n229, n230, n231, n232, n233, n234, n235, n236, n244, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U101 ( .A(n150), .B(n284), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n145), .B(n151), .CI(n100), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n166), .B(n153), .CI(n159), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  BUF_X2 U237 ( .A(n216), .Z(n333) );
  OAI21_X1 U238 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  OR2_X1 U239 ( .A1(n92), .A2(n95), .ZN(n274) );
  OR2_X1 U240 ( .A1(n172), .A2(n140), .ZN(n275) );
  XNOR2_X1 U241 ( .A(n308), .B(n276), .ZN(product[14]) );
  AND3_X1 U242 ( .A1(n305), .A2(n306), .A3(n307), .ZN(n276) );
  CLKBUF_X1 U243 ( .A(n236), .Z(n294) );
  NOR2_X1 U244 ( .A1(n92), .A2(n95), .ZN(n277) );
  NOR2_X1 U245 ( .A1(n92), .A2(n95), .ZN(n30) );
  OR2_X1 U246 ( .A1(n114), .A2(n117), .ZN(n278) );
  NOR2_X2 U247 ( .A1(n108), .A2(n113), .ZN(n44) );
  CLKBUF_X1 U248 ( .A(n333), .Z(n279) );
  CLKBUF_X1 U249 ( .A(n29), .Z(n280) );
  NAND2_X1 U250 ( .A1(n218), .A2(n226), .ZN(n281) );
  NAND2_X1 U251 ( .A1(n226), .A2(n218), .ZN(n222) );
  OAI21_X1 U252 ( .B1(n45), .B2(n41), .A(n42), .ZN(n40) );
  AND2_X1 U253 ( .A1(n118), .A2(n121), .ZN(n52) );
  BUF_X2 U254 ( .A(n233), .Z(n282) );
  CLKBUF_X1 U255 ( .A(n234), .Z(n283) );
  OAI22_X1 U256 ( .A1(n329), .A2(n192), .B1(n191), .B2(n297), .ZN(n284) );
  INV_X1 U257 ( .A(n126), .ZN(n285) );
  AND3_X1 U258 ( .A1(n311), .A2(n310), .A3(n309), .ZN(product[15]) );
  CLKBUF_X1 U259 ( .A(n39), .Z(n287) );
  CLKBUF_X1 U260 ( .A(n70), .Z(n288) );
  CLKBUF_X1 U261 ( .A(n47), .Z(n289) );
  INV_X1 U262 ( .A(n34), .ZN(n290) );
  CLKBUF_X1 U263 ( .A(n40), .Z(n291) );
  AOI21_X1 U264 ( .B1(n289), .B2(n287), .A(n291), .ZN(n292) );
  NAND2_X2 U265 ( .A1(n220), .A2(n244), .ZN(n293) );
  NAND2_X1 U266 ( .A1(n220), .A2(n244), .ZN(n224) );
  CLKBUF_X1 U267 ( .A(n235), .Z(n295) );
  INV_X1 U268 ( .A(n313), .ZN(n296) );
  INV_X1 U269 ( .A(n296), .ZN(n297) );
  INV_X1 U270 ( .A(n296), .ZN(n298) );
  NAND2_X2 U271 ( .A1(n217), .A2(n225), .ZN(n221) );
  NAND2_X1 U272 ( .A1(n236), .A2(n300), .ZN(n301) );
  NAND2_X1 U273 ( .A1(n299), .A2(n135), .ZN(n302) );
  NAND2_X1 U274 ( .A1(n301), .A2(n302), .ZN(n220) );
  INV_X1 U275 ( .A(n236), .ZN(n299) );
  INV_X1 U276 ( .A(n135), .ZN(n300) );
  INV_X1 U277 ( .A(n230), .ZN(n303) );
  XOR2_X1 U278 ( .A(n85), .B(n84), .Z(n304) );
  XOR2_X1 U279 ( .A(n304), .B(n288), .Z(product[13]) );
  NAND2_X1 U280 ( .A1(n85), .A2(n84), .ZN(n305) );
  NAND2_X1 U281 ( .A1(n85), .A2(n70), .ZN(n306) );
  NAND2_X1 U282 ( .A1(n70), .A2(n84), .ZN(n307) );
  NAND3_X1 U283 ( .A1(n306), .A2(n307), .A3(n305), .ZN(n14) );
  XOR2_X1 U284 ( .A(n141), .B(n83), .Z(n308) );
  NAND2_X1 U285 ( .A1(n141), .A2(n83), .ZN(n309) );
  NAND2_X1 U286 ( .A1(n14), .A2(n141), .ZN(n310) );
  NAND2_X1 U287 ( .A1(n14), .A2(n83), .ZN(n311) );
  XNOR2_X1 U288 ( .A(n236), .B(a[2]), .ZN(n313) );
  CLKBUF_X1 U289 ( .A(n20), .Z(n312) );
  XNOR2_X1 U290 ( .A(n236), .B(a[2]), .ZN(n227) );
  XNOR2_X1 U291 ( .A(n234), .B(a[6]), .ZN(n314) );
  INV_X1 U292 ( .A(n35), .ZN(n74) );
  XOR2_X1 U293 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U294 ( .A1(n274), .A2(n31), .ZN(n3) );
  AOI21_X1 U295 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XNOR2_X1 U296 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U297 ( .A1(n74), .A2(n290), .ZN(n4) );
  INV_X1 U298 ( .A(n36), .ZN(n34) );
  INV_X1 U299 ( .A(n26), .ZN(n24) );
  AOI21_X1 U300 ( .B1(n317), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U301 ( .A(n66), .ZN(n64) );
  NAND2_X1 U302 ( .A1(n318), .A2(n54), .ZN(n8) );
  NAND2_X1 U303 ( .A1(n320), .A2(n19), .ZN(n1) );
  XOR2_X1 U304 ( .A(n10), .B(n62), .Z(product[3]) );
  NAND2_X1 U305 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U306 ( .A(n60), .ZN(n80) );
  XOR2_X1 U307 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U308 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U309 ( .A(n56), .ZN(n79) );
  XOR2_X1 U310 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U311 ( .A1(n319), .A2(n26), .ZN(n2) );
  XOR2_X1 U312 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U313 ( .A1(n76), .A2(n45), .ZN(n6) );
  INV_X1 U314 ( .A(n44), .ZN(n76) );
  XNOR2_X1 U315 ( .A(n43), .B(n5), .ZN(product[8]) );
  OAI21_X1 U316 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U317 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U318 ( .A1(n317), .A2(n66), .ZN(n11) );
  OAI21_X1 U319 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  NAND2_X1 U320 ( .A1(n278), .A2(n49), .ZN(n7) );
  INV_X1 U321 ( .A(n19), .ZN(n17) );
  XNOR2_X1 U322 ( .A(n104), .B(n315), .ZN(n102) );
  XNOR2_X1 U323 ( .A(n106), .B(n109), .ZN(n315) );
  XNOR2_X1 U324 ( .A(n316), .B(n94), .ZN(n92) );
  XNOR2_X1 U325 ( .A(n97), .B(n144), .ZN(n316) );
  NOR2_X1 U326 ( .A1(n124), .A2(n139), .ZN(n60) );
  NAND2_X1 U327 ( .A1(n124), .A2(n139), .ZN(n61) );
  INV_X1 U328 ( .A(n69), .ZN(n67) );
  OR2_X1 U329 ( .A1(n171), .A2(n164), .ZN(n317) );
  NOR2_X1 U330 ( .A1(n122), .A2(n123), .ZN(n56) );
  OR2_X1 U331 ( .A1(n158), .A2(n146), .ZN(n105) );
  NOR2_X1 U332 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U333 ( .A(n83), .ZN(n84) );
  OR2_X1 U334 ( .A1(n118), .A2(n121), .ZN(n318) );
  OR2_X1 U335 ( .A1(n88), .A2(n91), .ZN(n319) );
  NAND2_X1 U336 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U337 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U338 ( .A1(n122), .A2(n123), .ZN(n57) );
  OR2_X1 U339 ( .A1(n87), .A2(n86), .ZN(n320) );
  NAND2_X1 U340 ( .A1(n118), .A2(n121), .ZN(n54) );
  OR2_X1 U341 ( .A1(n333), .A2(n231), .ZN(n199) );
  AND2_X1 U342 ( .A1(n333), .A2(n126), .ZN(n148) );
  AND2_X1 U343 ( .A1(n279), .A2(n129), .ZN(n156) );
  OR2_X1 U344 ( .A1(n333), .A2(n230), .ZN(n190) );
  INV_X1 U345 ( .A(n131), .ZN(n157) );
  INV_X1 U346 ( .A(n89), .ZN(n90) );
  INV_X1 U347 ( .A(n125), .ZN(n141) );
  INV_X1 U348 ( .A(n99), .ZN(n100) );
  OR2_X1 U349 ( .A1(n333), .A2(n229), .ZN(n181) );
  INV_X1 U350 ( .A(n128), .ZN(n149) );
  AND2_X1 U351 ( .A1(n333), .A2(n296), .ZN(n164) );
  AND2_X1 U352 ( .A1(n275), .A2(n69), .ZN(product[1]) );
  XNOR2_X1 U353 ( .A(n234), .B(a[6]), .ZN(n225) );
  OR2_X1 U354 ( .A1(n333), .A2(n232), .ZN(n208) );
  XNOR2_X1 U355 ( .A(n282), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U356 ( .A(n282), .B(b[4]), .ZN(n176) );
  XOR2_X1 U357 ( .A(n233), .B(a[6]), .Z(n217) );
  INV_X1 U358 ( .A(n135), .ZN(n244) );
  XNOR2_X1 U359 ( .A(n282), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U360 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U361 ( .A(n282), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U362 ( .A(n282), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U363 ( .A(n333), .B(n282), .ZN(n180) );
  INV_X1 U364 ( .A(n233), .ZN(n229) );
  AND2_X1 U365 ( .A1(n279), .A2(n135), .ZN(product[0]) );
  OAI22_X1 U366 ( .A1(n293), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  OAI22_X1 U367 ( .A1(n293), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U368 ( .A1(n293), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U369 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI22_X1 U370 ( .A1(n293), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U371 ( .A1(n293), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  INV_X1 U372 ( .A(n59), .ZN(n58) );
  NAND2_X1 U373 ( .A1(n104), .A2(n106), .ZN(n322) );
  NAND2_X1 U374 ( .A1(n104), .A2(n109), .ZN(n323) );
  NAND2_X1 U375 ( .A1(n106), .A2(n109), .ZN(n324) );
  NAND3_X1 U376 ( .A1(n322), .A2(n323), .A3(n324), .ZN(n101) );
  XNOR2_X1 U377 ( .A(n158), .B(n146), .ZN(n106) );
  INV_X1 U378 ( .A(n134), .ZN(n165) );
  NAND2_X1 U379 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI22_X1 U380 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U381 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  NOR2_X1 U382 ( .A1(n102), .A2(n107), .ZN(n325) );
  NOR2_X1 U383 ( .A1(n102), .A2(n107), .ZN(n41) );
  NAND2_X1 U384 ( .A1(n94), .A2(n97), .ZN(n326) );
  NAND2_X1 U385 ( .A1(n94), .A2(n144), .ZN(n327) );
  NAND2_X1 U386 ( .A1(n97), .A2(n144), .ZN(n328) );
  NAND3_X1 U387 ( .A1(n326), .A2(n327), .A3(n328), .ZN(n91) );
  NAND2_X1 U388 ( .A1(n219), .A2(n227), .ZN(n329) );
  NAND2_X1 U389 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U390 ( .A1(n219), .A2(n227), .ZN(n223) );
  AOI21_X1 U391 ( .B1(n318), .B2(n55), .A(n52), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n235), .B(a[4]), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n235), .B(a[4]), .ZN(n332) );
  AOI21_X1 U394 ( .B1(n318), .B2(n55), .A(n52), .ZN(n50) );
  XNOR2_X1 U395 ( .A(n235), .B(a[4]), .ZN(n226) );
  NAND2_X1 U396 ( .A1(n108), .A2(n113), .ZN(n45) );
  NAND2_X1 U397 ( .A1(n171), .A2(n164), .ZN(n66) );
  OAI22_X1 U398 ( .A1(n293), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  NAND2_X1 U399 ( .A1(n102), .A2(n107), .ZN(n42) );
  NAND2_X1 U400 ( .A1(n96), .A2(n101), .ZN(n36) );
  NAND2_X1 U401 ( .A1(n92), .A2(n95), .ZN(n31) );
  NAND2_X1 U402 ( .A1(n28), .A2(n319), .ZN(n21) );
  NOR2_X1 U403 ( .A1(n96), .A2(n101), .ZN(n35) );
  XNOR2_X1 U404 ( .A(n282), .B(b[7]), .ZN(n173) );
  OAI21_X1 U405 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  XNOR2_X1 U406 ( .A(n55), .B(n8), .ZN(product[5]) );
  OAI21_X1 U407 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  XNOR2_X1 U408 ( .A(n294), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U409 ( .A(n236), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U410 ( .A(n294), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U411 ( .A(n333), .B(n294), .ZN(n207) );
  XNOR2_X1 U412 ( .A(n236), .B(b[7]), .ZN(n200) );
  INV_X1 U413 ( .A(n236), .ZN(n232) );
  XNOR2_X1 U414 ( .A(n236), .B(b[1]), .ZN(n206) );
  XNOR2_X1 U415 ( .A(n294), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U416 ( .A(n236), .B(b[3]), .ZN(n204) );
  AOI21_X1 U417 ( .B1(n37), .B2(n28), .A(n280), .ZN(n27) );
  AOI21_X1 U418 ( .B1(n29), .B2(n319), .A(n24), .ZN(n22) );
  OAI21_X1 U419 ( .B1(n277), .B2(n36), .A(n31), .ZN(n29) );
  NOR2_X1 U420 ( .A1(n35), .A2(n30), .ZN(n28) );
  INV_X1 U421 ( .A(n289), .ZN(n46) );
  AOI21_X1 U422 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U423 ( .A1(n172), .A2(n140), .ZN(n69) );
  XOR2_X1 U424 ( .A(n7), .B(n330), .Z(product[6]) );
  OAI22_X1 U425 ( .A1(n182), .A2(n281), .B1(n182), .B2(n331), .ZN(n128) );
  OAI22_X1 U426 ( .A1(n281), .A2(n188), .B1(n187), .B2(n332), .ZN(n154) );
  OAI22_X1 U427 ( .A1(n281), .A2(n183), .B1(n182), .B2(n331), .ZN(n89) );
  OAI22_X1 U428 ( .A1(n281), .A2(n186), .B1(n185), .B2(n332), .ZN(n152) );
  OAI22_X1 U429 ( .A1(n187), .A2(n222), .B1(n186), .B2(n332), .ZN(n153) );
  OAI22_X1 U430 ( .A1(n281), .A2(n185), .B1(n184), .B2(n332), .ZN(n151) );
  OAI22_X1 U431 ( .A1(n281), .A2(n184), .B1(n183), .B2(n331), .ZN(n150) );
  INV_X1 U432 ( .A(n331), .ZN(n129) );
  XNOR2_X1 U433 ( .A(n235), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U434 ( .A(n235), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U435 ( .A(n235), .B(b[3]), .ZN(n195) );
  OAI22_X1 U436 ( .A1(n222), .A2(n230), .B1(n190), .B2(n332), .ZN(n138) );
  OAI22_X1 U437 ( .A1(n222), .A2(n189), .B1(n188), .B2(n331), .ZN(n155) );
  XNOR2_X1 U438 ( .A(n295), .B(b[2]), .ZN(n196) );
  INV_X1 U439 ( .A(n295), .ZN(n231) );
  XNOR2_X1 U440 ( .A(n235), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U441 ( .A(n235), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U442 ( .A(n333), .B(n295), .ZN(n198) );
  XNOR2_X1 U443 ( .A(n235), .B(b[1]), .ZN(n197) );
  XOR2_X1 U444 ( .A(n235), .B(a[2]), .Z(n219) );
  INV_X1 U445 ( .A(n325), .ZN(n75) );
  INV_X1 U446 ( .A(n15), .ZN(n70) );
  OAI22_X1 U447 ( .A1(n173), .A2(n221), .B1(n173), .B2(n285), .ZN(n125) );
  OAI22_X1 U448 ( .A1(n221), .A2(n174), .B1(n173), .B2(n285), .ZN(n83) );
  NOR2_X1 U449 ( .A1(n325), .A2(n44), .ZN(n39) );
  OAI22_X1 U450 ( .A1(n221), .A2(n175), .B1(n174), .B2(n285), .ZN(n142) );
  OAI22_X1 U451 ( .A1(n221), .A2(n176), .B1(n175), .B2(n285), .ZN(n143) );
  OAI22_X1 U452 ( .A1(n221), .A2(n177), .B1(n176), .B2(n285), .ZN(n144) );
  XNOR2_X1 U453 ( .A(n303), .B(b[7]), .ZN(n182) );
  OAI22_X1 U454 ( .A1(n221), .A2(n178), .B1(n177), .B2(n314), .ZN(n145) );
  INV_X1 U455 ( .A(n314), .ZN(n126) );
  OAI22_X1 U456 ( .A1(n221), .A2(n179), .B1(n178), .B2(n314), .ZN(n146) );
  XNOR2_X1 U457 ( .A(n283), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U458 ( .A(n283), .B(b[5]), .ZN(n184) );
  OAI22_X1 U459 ( .A1(n221), .A2(n229), .B1(n181), .B2(n314), .ZN(n137) );
  OAI22_X1 U460 ( .A1(n180), .A2(n221), .B1(n179), .B2(n314), .ZN(n147) );
  XNOR2_X1 U461 ( .A(n303), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U462 ( .A(n234), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U463 ( .A(n283), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U464 ( .A(n333), .B(n283), .ZN(n189) );
  INV_X1 U465 ( .A(n234), .ZN(n230) );
  XNOR2_X1 U466 ( .A(n234), .B(b[1]), .ZN(n188) );
  XOR2_X1 U467 ( .A(n234), .B(a[4]), .Z(n218) );
  XNOR2_X1 U468 ( .A(n312), .B(n1), .ZN(product[12]) );
  INV_X1 U469 ( .A(n292), .ZN(n37) );
  AOI21_X1 U470 ( .B1(n20), .B2(n320), .A(n17), .ZN(n15) );
  OAI22_X1 U471 ( .A1(n329), .A2(n193), .B1(n192), .B2(n297), .ZN(n158) );
  OAI22_X1 U472 ( .A1(n223), .A2(n195), .B1(n194), .B2(n297), .ZN(n160) );
  OAI22_X1 U473 ( .A1(n223), .A2(n194), .B1(n193), .B2(n227), .ZN(n159) );
  OAI22_X1 U474 ( .A1(n329), .A2(n196), .B1(n195), .B2(n298), .ZN(n161) );
  OAI22_X1 U475 ( .A1(n329), .A2(n231), .B1(n199), .B2(n297), .ZN(n139) );
  OAI22_X1 U476 ( .A1(n329), .A2(n197), .B1(n196), .B2(n298), .ZN(n162) );
  OAI22_X1 U477 ( .A1(n223), .A2(n192), .B1(n191), .B2(n298), .ZN(n99) );
  OAI22_X1 U478 ( .A1(n191), .A2(n329), .B1(n191), .B2(n297), .ZN(n131) );
  OAI22_X1 U479 ( .A1(n223), .A2(n198), .B1(n197), .B2(n297), .ZN(n163) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_8_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n54,
         n56, n57, n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  FA_X1 U6 ( .A(A[11]), .B(B[11]), .CI(n17), .CO(n16), .S(SUM[11]) );
  OR2_X1 U86 ( .A1(A[0]), .A2(B[0]), .ZN(n125) );
  AOI21_X1 U87 ( .B1(n137), .B2(n57), .A(n54), .ZN(n126) );
  AOI21_X1 U88 ( .B1(n137), .B2(n57), .A(n54), .ZN(n52) );
  AOI21_X1 U89 ( .B1(n33), .B2(n139), .A(n30), .ZN(n127) );
  CLKBUF_X1 U90 ( .A(n25), .Z(n128) );
  CLKBUF_X1 U91 ( .A(n41), .Z(n129) );
  CLKBUF_X1 U92 ( .A(n49), .Z(n130) );
  AOI21_X1 U93 ( .B1(n128), .B2(n140), .A(n22), .ZN(n131) );
  AOI21_X1 U94 ( .B1(n130), .B2(n136), .A(n46), .ZN(n132) );
  AOI21_X1 U95 ( .B1(n129), .B2(n138), .A(n38), .ZN(n133) );
  CLKBUF_X1 U96 ( .A(n33), .Z(n134) );
  INV_X1 U97 ( .A(n40), .ZN(n38) );
  INV_X1 U98 ( .A(n56), .ZN(n54) );
  AOI21_X1 U99 ( .B1(n25), .B2(n140), .A(n22), .ZN(n20) );
  INV_X1 U100 ( .A(n24), .ZN(n22) );
  AOI21_X1 U101 ( .B1(n33), .B2(n139), .A(n30), .ZN(n28) );
  INV_X1 U102 ( .A(n32), .ZN(n30) );
  AOI21_X1 U103 ( .B1(n49), .B2(n136), .A(n46), .ZN(n44) );
  INV_X1 U104 ( .A(n48), .ZN(n46) );
  NAND2_X1 U105 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U106 ( .A(n42), .ZN(n66) );
  NAND2_X1 U107 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U108 ( .A(n34), .ZN(n64) );
  NAND2_X1 U109 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U110 ( .A(n26), .ZN(n62) );
  NAND2_X1 U111 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U112 ( .A(n18), .ZN(n60) );
  NAND2_X1 U113 ( .A1(n136), .A2(n48), .ZN(n9) );
  NAND2_X1 U114 ( .A1(n138), .A2(n40), .ZN(n7) );
  XOR2_X1 U115 ( .A(n126), .B(n10), .Z(SUM[2]) );
  NAND2_X1 U116 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U117 ( .A(n50), .ZN(n68) );
  XNOR2_X1 U118 ( .A(n134), .B(n5), .ZN(SUM[7]) );
  NAND2_X1 U119 ( .A1(n139), .A2(n32), .ZN(n5) );
  XNOR2_X1 U120 ( .A(n128), .B(n3), .ZN(SUM[9]) );
  NAND2_X1 U121 ( .A1(n140), .A2(n24), .ZN(n3) );
  INV_X1 U122 ( .A(n59), .ZN(n57) );
  XNOR2_X1 U123 ( .A(n11), .B(n57), .ZN(SUM[1]) );
  NAND2_X1 U124 ( .A1(n137), .A2(n56), .ZN(n11) );
  XNOR2_X1 U125 ( .A(n13), .B(n135), .ZN(SUM[15]) );
  XNOR2_X1 U126 ( .A(B[15]), .B(A[15]), .ZN(n135) );
  OR2_X1 U127 ( .A1(A[3]), .A2(B[3]), .ZN(n136) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U129 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  NOR2_X1 U130 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U131 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U132 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  OR2_X1 U133 ( .A1(A[1]), .A2(B[1]), .ZN(n137) );
  NAND2_X1 U134 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U135 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U136 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U137 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  OR2_X1 U138 ( .A1(A[5]), .A2(B[5]), .ZN(n138) );
  OR2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(n139) );
  OR2_X1 U140 ( .A1(A[9]), .A2(B[9]), .ZN(n140) );
  NAND2_X1 U141 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  NAND2_X1 U142 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U143 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U144 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U145 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  AND2_X1 U146 ( .A1(n125), .A2(n59), .ZN(SUM[0]) );
  AOI21_X1 U147 ( .B1(n41), .B2(n138), .A(n38), .ZN(n36) );
  XNOR2_X1 U148 ( .A(n129), .B(n7), .ZN(SUM[5]) );
  XOR2_X1 U149 ( .A(n133), .B(n6), .Z(SUM[6]) );
  XOR2_X1 U150 ( .A(n132), .B(n8), .Z(SUM[4]) );
  OAI21_X1 U151 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  OAI21_X1 U152 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  NAND2_X1 U153 ( .A1(A[0]), .A2(B[0]), .ZN(n59) );
  XOR2_X1 U154 ( .A(n131), .B(n2), .Z(SUM[10]) );
  XNOR2_X1 U155 ( .A(n130), .B(n9), .ZN(SUM[3]) );
  XOR2_X1 U156 ( .A(n127), .B(n4), .Z(SUM[8]) );
  OAI21_X1 U157 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  NAND2_X1 U158 ( .A1(A[1]), .A2(B[1]), .ZN(n56) );
  OAI21_X1 U159 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X1 U160 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
endmodule


module add_layer_WIDTH16_8 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_8_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n56,
         n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  FA_X1 U6 ( .A(A[11]), .B(B[11]), .CI(n17), .CO(n16), .S(SUM[11]) );
  AND2_X1 U86 ( .A1(A[1]), .A2(B[1]), .ZN(n128) );
  INV_X1 U87 ( .A(n127), .ZN(n59) );
  INV_X1 U88 ( .A(n128), .ZN(n56) );
  OR2_X1 U89 ( .A1(A[0]), .A2(B[0]), .ZN(n125) );
  AOI21_X1 U90 ( .B1(n49), .B2(n139), .A(n46), .ZN(n126) );
  AND2_X2 U91 ( .A1(A[0]), .A2(B[0]), .ZN(n127) );
  OR2_X2 U92 ( .A1(A[1]), .A2(B[1]), .ZN(n136) );
  AOI21_X1 U93 ( .B1(n49), .B2(n139), .A(n46), .ZN(n44) );
  CLKBUF_X1 U94 ( .A(n25), .Z(n129) );
  AOI21_X1 U95 ( .B1(n136), .B2(n127), .A(n128), .ZN(n130) );
  CLKBUF_X1 U96 ( .A(n41), .Z(n131) );
  CLKBUF_X1 U97 ( .A(n33), .Z(n132) );
  AOI21_X1 U98 ( .B1(n131), .B2(n140), .A(n38), .ZN(n133) );
  AOI21_X1 U99 ( .B1(n41), .B2(n140), .A(n38), .ZN(n36) );
  AOI21_X1 U100 ( .B1(n129), .B2(n141), .A(n22), .ZN(n134) );
  AOI21_X1 U101 ( .B1(n132), .B2(n138), .A(n30), .ZN(n135) );
  INV_X1 U102 ( .A(n32), .ZN(n30) );
  INV_X1 U103 ( .A(n48), .ZN(n46) );
  INV_X1 U104 ( .A(n40), .ZN(n38) );
  AOI21_X1 U105 ( .B1(n25), .B2(n141), .A(n22), .ZN(n20) );
  INV_X1 U106 ( .A(n24), .ZN(n22) );
  NAND2_X1 U107 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U108 ( .A(n42), .ZN(n66) );
  NAND2_X1 U109 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U110 ( .A(n34), .ZN(n64) );
  NAND2_X1 U111 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U112 ( .A(n26), .ZN(n62) );
  AOI21_X1 U113 ( .B1(n136), .B2(n127), .A(n128), .ZN(n52) );
  NAND2_X1 U114 ( .A1(n140), .A2(n40), .ZN(n7) );
  NAND2_X1 U115 ( .A1(n138), .A2(n32), .ZN(n5) );
  NAND2_X1 U116 ( .A1(n139), .A2(n48), .ZN(n9) );
  XOR2_X1 U117 ( .A(n134), .B(n2), .Z(SUM[10]) );
  NAND2_X1 U118 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U119 ( .A(n18), .ZN(n60) );
  XNOR2_X1 U120 ( .A(n129), .B(n3), .ZN(SUM[9]) );
  NAND2_X1 U121 ( .A1(n141), .A2(n24), .ZN(n3) );
  XNOR2_X1 U122 ( .A(n11), .B(n127), .ZN(SUM[1]) );
  NAND2_X1 U123 ( .A1(n136), .A2(n56), .ZN(n11) );
  NAND2_X1 U124 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U125 ( .A(n50), .ZN(n68) );
  XNOR2_X1 U126 ( .A(n13), .B(n137), .ZN(SUM[15]) );
  XNOR2_X1 U127 ( .A(B[15]), .B(A[15]), .ZN(n137) );
  NOR2_X1 U128 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U129 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U130 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U131 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  NOR2_X1 U132 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U133 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U134 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U135 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U136 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  OR2_X1 U137 ( .A1(A[7]), .A2(B[7]), .ZN(n138) );
  OR2_X1 U138 ( .A1(A[3]), .A2(B[3]), .ZN(n139) );
  OR2_X1 U139 ( .A1(A[5]), .A2(B[5]), .ZN(n140) );
  OR2_X1 U140 ( .A1(A[9]), .A2(B[9]), .ZN(n141) );
  NAND2_X1 U141 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  NAND2_X1 U142 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U143 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U144 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U145 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  AND2_X1 U146 ( .A1(n125), .A2(n59), .ZN(SUM[0]) );
  XNOR2_X1 U147 ( .A(n131), .B(n7), .ZN(SUM[5]) );
  XNOR2_X1 U148 ( .A(n49), .B(n9), .ZN(SUM[3]) );
  XOR2_X1 U149 ( .A(n126), .B(n8), .Z(SUM[4]) );
  OAI21_X1 U150 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  XNOR2_X1 U151 ( .A(n132), .B(n5), .ZN(SUM[7]) );
  XOR2_X1 U152 ( .A(n130), .B(n10), .Z(SUM[2]) );
  AOI21_X1 U153 ( .B1(n33), .B2(n138), .A(n30), .ZN(n28) );
  OAI21_X1 U154 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X1 U155 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  XOR2_X1 U156 ( .A(n133), .B(n6), .Z(SUM[6]) );
  OAI21_X1 U157 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U158 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U159 ( .A(n135), .B(n4), .Z(SUM[8]) );
endmodule


module add_layer_WIDTH16_7 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_7_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n21,
         n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37, n38, n39,
         n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55, n56, n57,
         n61, n64, n65, n67, n69, n71, n73, n75, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n173;

  NAND2_X1 U94 ( .A1(A[13]), .A2(B[13]), .ZN(n150) );
  OR2_X1 U95 ( .A1(A[0]), .A2(B[0]), .ZN(n132) );
  OAI21_X1 U96 ( .B1(n136), .B2(n137), .A(n21), .ZN(n133) );
  CLKBUF_X1 U97 ( .A(n46), .Z(n134) );
  CLKBUF_X1 U98 ( .A(n49), .Z(n135) );
  AOI21_X1 U99 ( .B1(n54), .B2(n168), .A(n51), .ZN(n49) );
  OAI21_X1 U100 ( .B1(n136), .B2(n137), .A(n21), .ZN(n65) );
  INV_X1 U101 ( .A(n170), .ZN(n136) );
  INV_X1 U102 ( .A(n22), .ZN(n137) );
  AOI21_X1 U103 ( .B1(n134), .B2(n169), .A(n43), .ZN(n138) );
  AOI21_X1 U104 ( .B1(n46), .B2(n169), .A(n43), .ZN(n41) );
  CLKBUF_X1 U105 ( .A(n54), .Z(n139) );
  CLKBUF_X1 U106 ( .A(n133), .Z(n140) );
  XOR2_X1 U107 ( .A(A[12]), .B(B[12]), .Z(n141) );
  XOR2_X1 U108 ( .A(n140), .B(n141), .Z(SUM[12]) );
  NAND2_X1 U109 ( .A1(n133), .A2(A[12]), .ZN(n142) );
  NAND2_X1 U110 ( .A1(n65), .A2(B[12]), .ZN(n143) );
  NAND2_X1 U111 ( .A1(A[12]), .A2(B[12]), .ZN(n144) );
  NAND3_X1 U112 ( .A1(n142), .A2(n143), .A3(n144), .ZN(n16) );
  CLKBUF_X1 U113 ( .A(n151), .Z(n145) );
  NAND3_X1 U114 ( .A1(n145), .A2(n150), .A3(n152), .ZN(n146) );
  CLKBUF_X1 U115 ( .A(n16), .Z(n147) );
  NAND3_X1 U116 ( .A1(n152), .A2(n151), .A3(n150), .ZN(n148) );
  XOR2_X1 U117 ( .A(A[13]), .B(B[13]), .Z(n149) );
  XOR2_X1 U118 ( .A(n149), .B(n147), .Z(SUM[13]) );
  NAND2_X1 U119 ( .A1(n16), .A2(A[13]), .ZN(n151) );
  NAND2_X1 U120 ( .A1(n16), .A2(B[13]), .ZN(n152) );
  NAND3_X1 U121 ( .A1(n152), .A2(n151), .A3(n150), .ZN(n15) );
  XOR2_X1 U122 ( .A(A[14]), .B(B[14]), .Z(n153) );
  XOR2_X1 U123 ( .A(n153), .B(n146), .Z(SUM[14]) );
  NAND2_X1 U124 ( .A1(A[14]), .A2(B[14]), .ZN(n154) );
  NAND2_X1 U125 ( .A1(n148), .A2(A[14]), .ZN(n155) );
  NAND2_X1 U126 ( .A1(n15), .A2(B[14]), .ZN(n156) );
  NAND3_X1 U127 ( .A1(n156), .A2(n155), .A3(n154), .ZN(n14) );
  OR2_X1 U128 ( .A1(A[1]), .A2(B[1]), .ZN(n157) );
  INV_X1 U129 ( .A(n61), .ZN(n158) );
  OR2_X1 U130 ( .A1(A[1]), .A2(B[1]), .ZN(n171) );
  AND2_X1 U131 ( .A1(A[1]), .A2(B[1]), .ZN(n163) );
  INV_X1 U132 ( .A(n163), .ZN(n61) );
  AND2_X1 U133 ( .A1(A[0]), .A2(B[0]), .ZN(n159) );
  CLKBUF_X1 U134 ( .A(n22), .Z(n160) );
  CLKBUF_X1 U135 ( .A(n30), .Z(n161) );
  CLKBUF_X1 U136 ( .A(n38), .Z(n162) );
  AOI21_X1 U137 ( .B1(n38), .B2(n167), .A(n35), .ZN(n164) );
  AOI21_X1 U138 ( .B1(n171), .B2(n159), .A(n163), .ZN(n165) );
  INV_X1 U139 ( .A(n53), .ZN(n51) );
  INV_X1 U140 ( .A(n45), .ZN(n43) );
  INV_X1 U141 ( .A(n37), .ZN(n35) );
  NAND2_X1 U142 ( .A1(n73), .A2(n48), .ZN(n9) );
  INV_X1 U143 ( .A(n47), .ZN(n73) );
  NAND2_X1 U144 ( .A1(n71), .A2(n40), .ZN(n7) );
  INV_X1 U145 ( .A(n39), .ZN(n71) );
  NAND2_X1 U146 ( .A1(n168), .A2(n53), .ZN(n10) );
  NAND2_X1 U147 ( .A1(n169), .A2(n45), .ZN(n8) );
  NAND2_X1 U148 ( .A1(n167), .A2(n37), .ZN(n6) );
  NAND2_X1 U149 ( .A1(n166), .A2(n29), .ZN(n4) );
  NAND2_X1 U150 ( .A1(n157), .A2(n61), .ZN(n12) );
  INV_X1 U151 ( .A(n29), .ZN(n27) );
  NAND2_X1 U152 ( .A1(n170), .A2(n21), .ZN(n2) );
  NAND2_X1 U153 ( .A1(n69), .A2(n32), .ZN(n5) );
  INV_X1 U154 ( .A(n31), .ZN(n69) );
  NAND2_X1 U155 ( .A1(n67), .A2(n24), .ZN(n3) );
  INV_X1 U156 ( .A(n23), .ZN(n67) );
  NAND2_X1 U157 ( .A1(n75), .A2(n56), .ZN(n11) );
  INV_X1 U158 ( .A(n55), .ZN(n75) );
  XOR2_X1 U159 ( .A(B[15]), .B(A[15]), .Z(n1) );
  OR2_X1 U160 ( .A1(A[9]), .A2(B[9]), .ZN(n166) );
  NOR2_X1 U161 ( .A1(A[6]), .A2(B[6]), .ZN(n39) );
  NOR2_X1 U162 ( .A1(A[8]), .A2(B[8]), .ZN(n31) );
  NOR2_X1 U163 ( .A1(A[2]), .A2(B[2]), .ZN(n55) );
  NOR2_X1 U164 ( .A1(A[4]), .A2(B[4]), .ZN(n47) );
  NOR2_X1 U165 ( .A1(A[10]), .A2(B[10]), .ZN(n23) );
  NAND2_X1 U166 ( .A1(A[9]), .A2(B[9]), .ZN(n29) );
  NAND2_X1 U167 ( .A1(A[7]), .A2(B[7]), .ZN(n37) );
  NAND2_X1 U168 ( .A1(A[3]), .A2(B[3]), .ZN(n53) );
  NAND2_X1 U169 ( .A1(A[5]), .A2(B[5]), .ZN(n45) );
  NAND2_X1 U170 ( .A1(A[11]), .A2(B[11]), .ZN(n21) );
  OR2_X1 U171 ( .A1(A[7]), .A2(B[7]), .ZN(n167) );
  OR2_X1 U172 ( .A1(A[3]), .A2(B[3]), .ZN(n168) );
  OR2_X1 U173 ( .A1(A[5]), .A2(B[5]), .ZN(n169) );
  OR2_X1 U174 ( .A1(A[11]), .A2(B[11]), .ZN(n170) );
  NAND2_X1 U175 ( .A1(A[6]), .A2(B[6]), .ZN(n40) );
  NAND2_X1 U176 ( .A1(A[8]), .A2(B[8]), .ZN(n32) );
  NAND2_X1 U177 ( .A1(A[2]), .A2(B[2]), .ZN(n56) );
  NAND2_X1 U178 ( .A1(A[4]), .A2(B[4]), .ZN(n48) );
  NAND2_X1 U179 ( .A1(A[10]), .A2(B[10]), .ZN(n24) );
  AND2_X1 U180 ( .A1(n132), .A2(n64), .ZN(SUM[0]) );
  XNOR2_X1 U181 ( .A(n134), .B(n8), .ZN(SUM[5]) );
  XNOR2_X1 U182 ( .A(n139), .B(n10), .ZN(SUM[3]) );
  XNOR2_X1 U183 ( .A(n12), .B(n159), .ZN(SUM[1]) );
  XOR2_X1 U184 ( .A(n135), .B(n9), .Z(SUM[4]) );
  XOR2_X1 U185 ( .A(n57), .B(n11), .Z(SUM[2]) );
  OAI21_X1 U186 ( .B1(n165), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U187 ( .B1(n157), .B2(n159), .A(n158), .ZN(n57) );
  AOI21_X1 U188 ( .B1(n162), .B2(n167), .A(n35), .ZN(n33) );
  OAI21_X1 U189 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U190 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  AOI21_X1 U191 ( .B1(n161), .B2(n166), .A(n27), .ZN(n173) );
  XOR2_X1 U192 ( .A(n14), .B(n1), .Z(SUM[15]) );
  NAND2_X1 U193 ( .A1(A[0]), .A2(B[0]), .ZN(n64) );
  XNOR2_X1 U194 ( .A(n161), .B(n4), .ZN(SUM[9]) );
  XOR2_X1 U195 ( .A(n33), .B(n5), .Z(SUM[8]) );
  AOI21_X1 U196 ( .B1(n30), .B2(n166), .A(n27), .ZN(n25) );
  OAI21_X1 U197 ( .B1(n164), .B2(n31), .A(n32), .ZN(n30) );
  XNOR2_X1 U198 ( .A(n162), .B(n6), .ZN(SUM[7]) );
  XOR2_X1 U199 ( .A(n173), .B(n3), .Z(SUM[10]) );
  XNOR2_X1 U200 ( .A(n160), .B(n2), .ZN(SUM[11]) );
  OAI21_X1 U201 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
  XOR2_X1 U202 ( .A(n138), .B(n7), .Z(SUM[6]) );
endmodule


module add_layer_WIDTH16_2 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_2_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_2 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_2 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_2 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_8 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_7 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_2 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_2 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8 \genblk1[0].mult  ( .clk(clk), .ia(
        {\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7 \genblk1[1].mult  ( .clk(clk), .ia(
        {\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6 \genblk1[2].mult  ( .clk(clk), .ia(
        {\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5 \genblk1[3].mult  ( .clk(clk), .ia(
        {\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_2 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n73,
         n74, n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n128, n129, n131, n132, n134, n135, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n229, n230, n231, n232, n233, n234, n235, n236,
         n244, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n324, n325, n326, n327, n328, n329,
         n330;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n150), .B(n302), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n145), .B(n100), .CI(n151), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n159), .B(n166), .CI(n153), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  FA_X1 U114 ( .A(n161), .B(n168), .CI(n120), .CO(n117), .S(n118) );
  HA_X1 U115 ( .A(n138), .B(n155), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n170), .B(n163), .CO(n123), .S(n124) );
  BUF_X2 U237 ( .A(n216), .Z(n330) );
  CLKBUF_X1 U238 ( .A(n35), .Z(n274) );
  AND2_X1 U239 ( .A1(n118), .A2(n121), .ZN(n277) );
  OR2_X1 U240 ( .A1(n88), .A2(n91), .ZN(n320) );
  INV_X1 U241 ( .A(n277), .ZN(n54) );
  OR2_X1 U242 ( .A1(n172), .A2(n140), .ZN(n275) );
  XNOR2_X1 U243 ( .A(n329), .B(b[7]), .ZN(n276) );
  CLKBUF_X3 U244 ( .A(n236), .Z(n329) );
  CLKBUF_X1 U245 ( .A(n36), .Z(n278) );
  NAND3_X1 U246 ( .A1(n309), .A2(n308), .A3(n307), .ZN(n279) );
  NOR2_X1 U247 ( .A1(n92), .A2(n95), .ZN(n280) );
  NOR2_X1 U248 ( .A1(n92), .A2(n95), .ZN(n30) );
  XNOR2_X1 U249 ( .A(n104), .B(n281), .ZN(n102) );
  XNOR2_X1 U250 ( .A(n109), .B(n106), .ZN(n281) );
  CLKBUF_X1 U251 ( .A(n325), .Z(n282) );
  NAND2_X1 U252 ( .A1(n14), .A2(n83), .ZN(n312) );
  NAND3_X1 U253 ( .A1(n309), .A2(n308), .A3(n307), .ZN(n14) );
  XOR2_X1 U254 ( .A(n234), .B(a[4]), .Z(n283) );
  CLKBUF_X1 U255 ( .A(n234), .Z(n284) );
  CLKBUF_X1 U256 ( .A(n235), .Z(n285) );
  XNOR2_X1 U257 ( .A(n235), .B(a[4]), .ZN(n286) );
  INV_X1 U258 ( .A(n73), .ZN(n287) );
  OAI21_X1 U259 ( .B1(n287), .B2(n278), .A(n31), .ZN(n288) );
  XOR2_X1 U260 ( .A(n235), .B(a[2]), .Z(n289) );
  BUF_X1 U261 ( .A(n226), .Z(n324) );
  AOI21_X1 U262 ( .B1(n319), .B2(n55), .A(n277), .ZN(n290) );
  AOI21_X1 U263 ( .B1(n319), .B2(n55), .A(n277), .ZN(n50) );
  CLKBUF_X1 U264 ( .A(n70), .Z(n291) );
  CLKBUF_X1 U265 ( .A(n28), .Z(n292) );
  XNOR2_X1 U266 ( .A(n234), .B(a[6]), .ZN(n293) );
  XNOR2_X1 U267 ( .A(n234), .B(a[6]), .ZN(n225) );
  BUF_X1 U268 ( .A(n326), .Z(n294) );
  XNOR2_X1 U269 ( .A(n295), .B(n301), .ZN(product[14]) );
  XNOR2_X1 U270 ( .A(n141), .B(n83), .ZN(n295) );
  BUF_X1 U271 ( .A(n225), .Z(n318) );
  NAND2_X1 U272 ( .A1(n104), .A2(n109), .ZN(n296) );
  NAND2_X1 U273 ( .A1(n104), .A2(n106), .ZN(n297) );
  NAND2_X1 U274 ( .A1(n109), .A2(n106), .ZN(n298) );
  NAND3_X1 U275 ( .A1(n296), .A2(n297), .A3(n298), .ZN(n101) );
  CLKBUF_X1 U276 ( .A(n40), .Z(n299) );
  CLKBUF_X1 U277 ( .A(n234), .Z(n300) );
  NAND3_X1 U278 ( .A1(n307), .A2(n308), .A3(n309), .ZN(n301) );
  OAI22_X1 U279 ( .A1(n223), .A2(n192), .B1(n191), .B2(n304), .ZN(n302) );
  BUF_X2 U280 ( .A(n227), .Z(n303) );
  BUF_X1 U281 ( .A(n227), .Z(n304) );
  XNOR2_X1 U282 ( .A(n236), .B(a[2]), .ZN(n227) );
  AND3_X1 U283 ( .A1(n310), .A2(n311), .A3(n312), .ZN(product[15]) );
  NAND2_X1 U284 ( .A1(n108), .A2(n113), .ZN(n45) );
  NAND2_X1 U285 ( .A1(n96), .A2(n101), .ZN(n36) );
  XOR2_X1 U286 ( .A(n85), .B(n84), .Z(n306) );
  XOR2_X1 U287 ( .A(n306), .B(n291), .Z(product[13]) );
  NAND2_X1 U288 ( .A1(n85), .A2(n84), .ZN(n307) );
  NAND2_X1 U289 ( .A1(n85), .A2(n70), .ZN(n308) );
  NAND2_X1 U290 ( .A1(n84), .A2(n70), .ZN(n309) );
  NAND2_X1 U291 ( .A1(n141), .A2(n83), .ZN(n310) );
  NAND2_X1 U292 ( .A1(n279), .A2(n141), .ZN(n311) );
  CLKBUF_X1 U293 ( .A(n20), .Z(n313) );
  CLKBUF_X1 U294 ( .A(n233), .Z(n314) );
  OAI21_X1 U295 ( .B1(n48), .B2(n290), .A(n49), .ZN(n315) );
  NOR2_X1 U296 ( .A1(n102), .A2(n107), .ZN(n316) );
  AOI21_X1 U297 ( .B1(n39), .B2(n315), .A(n299), .ZN(n317) );
  NOR2_X1 U298 ( .A1(n108), .A2(n113), .ZN(n44) );
  INV_X2 U299 ( .A(n135), .ZN(n244) );
  INV_X1 U300 ( .A(n274), .ZN(n74) );
  XNOR2_X1 U301 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U302 ( .A1(n74), .A2(n278), .ZN(n4) );
  INV_X1 U303 ( .A(n278), .ZN(n34) );
  AOI21_X1 U304 ( .B1(n321), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U305 ( .A(n26), .ZN(n24) );
  NAND2_X1 U306 ( .A1(n319), .A2(n54), .ZN(n8) );
  NAND2_X1 U307 ( .A1(n322), .A2(n19), .ZN(n1) );
  XOR2_X1 U308 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U309 ( .A1(n73), .A2(n31), .ZN(n3) );
  AOI21_X1 U310 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U311 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U312 ( .A1(n76), .A2(n45), .ZN(n6) );
  INV_X1 U313 ( .A(n44), .ZN(n76) );
  XOR2_X1 U314 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U315 ( .A1(n320), .A2(n26), .ZN(n2) );
  NOR2_X1 U316 ( .A1(n96), .A2(n101), .ZN(n35) );
  NOR2_X1 U317 ( .A1(n35), .A2(n280), .ZN(n28) );
  XNOR2_X1 U318 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U319 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U320 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U321 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U322 ( .A1(n321), .A2(n66), .ZN(n11) );
  NAND2_X1 U323 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U324 ( .A(n48), .ZN(n77) );
  INV_X1 U325 ( .A(n19), .ZN(n17) );
  OR2_X1 U326 ( .A1(n158), .A2(n146), .ZN(n105) );
  OAI21_X1 U327 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  OR2_X1 U328 ( .A1(n118), .A2(n121), .ZN(n319) );
  XOR2_X1 U329 ( .A(n10), .B(n62), .Z(product[3]) );
  NAND2_X1 U330 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U331 ( .A(n60), .ZN(n80) );
  XOR2_X1 U332 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U333 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U334 ( .A(n56), .ZN(n79) );
  XNOR2_X1 U335 ( .A(n158), .B(n146), .ZN(n106) );
  NOR2_X1 U336 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U337 ( .A(n83), .ZN(n84) );
  OAI21_X1 U338 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  OR2_X1 U339 ( .A1(n171), .A2(n164), .ZN(n321) );
  NAND2_X1 U340 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U341 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U342 ( .A1(n114), .A2(n117), .ZN(n49) );
  OR2_X1 U343 ( .A1(n87), .A2(n86), .ZN(n322) );
  INV_X1 U344 ( .A(n131), .ZN(n157) );
  INV_X1 U345 ( .A(n128), .ZN(n149) );
  INV_X1 U346 ( .A(n89), .ZN(n90) );
  OAI22_X1 U347 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  AND2_X1 U348 ( .A1(n330), .A2(n129), .ZN(n156) );
  OAI22_X1 U349 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  AND2_X1 U350 ( .A1(n330), .A2(n126), .ZN(n148) );
  OAI22_X1 U351 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OR2_X1 U352 ( .A1(n330), .A2(n230), .ZN(n190) );
  OAI22_X1 U353 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  NOR2_X1 U354 ( .A1(n124), .A2(n139), .ZN(n60) );
  NOR2_X1 U355 ( .A1(n122), .A2(n123), .ZN(n56) );
  INV_X1 U356 ( .A(n125), .ZN(n141) );
  NAND2_X1 U357 ( .A1(n122), .A2(n123), .ZN(n57) );
  AND2_X1 U358 ( .A1(n330), .A2(n132), .ZN(n164) );
  OR2_X1 U359 ( .A1(n330), .A2(n229), .ZN(n181) );
  AND2_X1 U360 ( .A1(n275), .A2(n69), .ZN(product[1]) );
  OR2_X1 U361 ( .A1(n330), .A2(n232), .ZN(n208) );
  XNOR2_X1 U362 ( .A(n330), .B(n233), .ZN(n180) );
  XNOR2_X1 U363 ( .A(n314), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U364 ( .A(n314), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U365 ( .A(n233), .B(b[2]), .ZN(n178) );
  INV_X1 U366 ( .A(n233), .ZN(n229) );
  AND2_X1 U367 ( .A1(n330), .A2(n135), .ZN(product[0]) );
  XNOR2_X1 U368 ( .A(n235), .B(a[4]), .ZN(n226) );
  NAND2_X1 U369 ( .A1(n171), .A2(n164), .ZN(n66) );
  NAND2_X1 U370 ( .A1(n124), .A2(n139), .ZN(n61) );
  NAND2_X1 U371 ( .A1(n172), .A2(n140), .ZN(n69) );
  NAND2_X1 U372 ( .A1(n217), .A2(n225), .ZN(n325) );
  NAND2_X1 U373 ( .A1(n217), .A2(n293), .ZN(n221) );
  XNOR2_X1 U374 ( .A(n314), .B(b[6]), .ZN(n174) );
  OR2_X1 U375 ( .A1(n330), .A2(n231), .ZN(n199) );
  NAND2_X1 U376 ( .A1(n219), .A2(n227), .ZN(n223) );
  NAND2_X1 U377 ( .A1(n289), .A2(n227), .ZN(n328) );
  NAND2_X1 U378 ( .A1(n226), .A2(n218), .ZN(n222) );
  NAND2_X1 U379 ( .A1(n283), .A2(n286), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n314), .B(b[7]), .ZN(n173) );
  XOR2_X1 U381 ( .A(n233), .B(a[6]), .Z(n217) );
  CLKBUF_X1 U382 ( .A(n235), .Z(n327) );
  AOI21_X1 U383 ( .B1(n37), .B2(n292), .A(n288), .ZN(n27) );
  INV_X1 U384 ( .A(n99), .ZN(n100) );
  XNOR2_X1 U385 ( .A(n8), .B(n55), .ZN(product[5]) );
  NAND2_X1 U386 ( .A1(n102), .A2(n107), .ZN(n42) );
  OAI22_X1 U387 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  INV_X1 U388 ( .A(n134), .ZN(n165) );
  OAI22_X1 U389 ( .A1(n276), .A2(n224), .B1(n276), .B2(n244), .ZN(n134) );
  OAI22_X1 U390 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  INV_X1 U391 ( .A(n59), .ZN(n58) );
  INV_X1 U392 ( .A(n66), .ZN(n64) );
  INV_X1 U393 ( .A(n69), .ZN(n67) );
  OAI22_X1 U394 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  NAND2_X2 U395 ( .A1(n220), .A2(n244), .ZN(n224) );
  XNOR2_X1 U396 ( .A(n300), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U397 ( .A(n234), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U398 ( .A(n284), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U399 ( .A(n300), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U400 ( .A(n234), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U401 ( .A(n330), .B(n284), .ZN(n189) );
  INV_X1 U402 ( .A(n234), .ZN(n230) );
  XOR2_X1 U403 ( .A(n234), .B(a[4]), .Z(n218) );
  INV_X1 U404 ( .A(n280), .ZN(n73) );
  OAI21_X1 U405 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  NAND2_X1 U406 ( .A1(n92), .A2(n95), .ZN(n31) );
  INV_X1 U407 ( .A(n316), .ZN(n75) );
  NOR2_X1 U408 ( .A1(n316), .A2(n44), .ZN(n39) );
  NOR2_X1 U409 ( .A1(n102), .A2(n107), .ZN(n41) );
  XNOR2_X1 U410 ( .A(n233), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U411 ( .A(n284), .B(b[3]), .ZN(n186) );
  NAND2_X1 U412 ( .A1(n28), .A2(n320), .ZN(n21) );
  OAI22_X1 U413 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI21_X1 U414 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U415 ( .B1(n29), .B2(n320), .A(n24), .ZN(n22) );
  OAI21_X1 U416 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  XNOR2_X1 U417 ( .A(n234), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U418 ( .A(n233), .B(b[1]), .ZN(n179) );
  XOR2_X1 U419 ( .A(n7), .B(n290), .Z(product[6]) );
  INV_X1 U420 ( .A(n315), .ZN(n46) );
  AOI21_X1 U421 ( .B1(n39), .B2(n47), .A(n40), .ZN(n38) );
  OAI21_X1 U422 ( .B1(n48), .B2(n50), .A(n49), .ZN(n47) );
  OAI22_X1 U423 ( .A1(n182), .A2(n294), .B1(n182), .B2(n324), .ZN(n128) );
  OAI22_X1 U424 ( .A1(n326), .A2(n183), .B1(n182), .B2(n324), .ZN(n89) );
  OAI22_X1 U425 ( .A1(n294), .A2(n188), .B1(n187), .B2(n286), .ZN(n154) );
  OAI22_X1 U426 ( .A1(n326), .A2(n185), .B1(n184), .B2(n286), .ZN(n151) );
  OAI22_X1 U427 ( .A1(n222), .A2(n187), .B1(n186), .B2(n286), .ZN(n153) );
  OAI22_X1 U428 ( .A1(n222), .A2(n184), .B1(n183), .B2(n286), .ZN(n150) );
  OAI22_X1 U429 ( .A1(n222), .A2(n186), .B1(n185), .B2(n324), .ZN(n152) );
  INV_X1 U430 ( .A(n324), .ZN(n129) );
  XNOR2_X1 U431 ( .A(n235), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U432 ( .A(n235), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U433 ( .A(n327), .B(b[3]), .ZN(n195) );
  OAI22_X1 U434 ( .A1(n222), .A2(n230), .B1(n190), .B2(n286), .ZN(n138) );
  OAI22_X1 U435 ( .A1(n222), .A2(n189), .B1(n188), .B2(n324), .ZN(n155) );
  XNOR2_X1 U436 ( .A(n327), .B(b[2]), .ZN(n196) );
  INV_X1 U437 ( .A(n285), .ZN(n231) );
  XNOR2_X1 U438 ( .A(n235), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U439 ( .A(n235), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U440 ( .A(n330), .B(n285), .ZN(n198) );
  XNOR2_X1 U441 ( .A(n285), .B(b[1]), .ZN(n197) );
  XOR2_X1 U442 ( .A(n235), .B(a[2]), .Z(n219) );
  INV_X1 U443 ( .A(n15), .ZN(n70) );
  OAI22_X1 U444 ( .A1(n173), .A2(n282), .B1(n173), .B2(n318), .ZN(n125) );
  OAI22_X1 U445 ( .A1(n282), .A2(n174), .B1(n173), .B2(n318), .ZN(n83) );
  OAI22_X1 U446 ( .A1(n282), .A2(n175), .B1(n174), .B2(n318), .ZN(n142) );
  OAI22_X1 U447 ( .A1(n282), .A2(n176), .B1(n175), .B2(n318), .ZN(n143) );
  OAI22_X1 U448 ( .A1(n325), .A2(n177), .B1(n176), .B2(n318), .ZN(n144) );
  OAI22_X1 U449 ( .A1(n325), .A2(n179), .B1(n178), .B2(n318), .ZN(n146) );
  OAI22_X1 U450 ( .A1(n325), .A2(n178), .B1(n177), .B2(n318), .ZN(n145) );
  INV_X1 U451 ( .A(n293), .ZN(n126) );
  OAI22_X1 U452 ( .A1(n221), .A2(n229), .B1(n181), .B2(n293), .ZN(n137) );
  OAI22_X1 U453 ( .A1(n221), .A2(n180), .B1(n179), .B2(n293), .ZN(n147) );
  XNOR2_X1 U454 ( .A(n313), .B(n1), .ZN(product[12]) );
  INV_X1 U455 ( .A(n317), .ZN(n37) );
  AOI21_X1 U456 ( .B1(n20), .B2(n322), .A(n17), .ZN(n15) );
  OAI22_X1 U457 ( .A1(n328), .A2(n193), .B1(n192), .B2(n304), .ZN(n158) );
  OAI22_X1 U458 ( .A1(n328), .A2(n195), .B1(n194), .B2(n303), .ZN(n160) );
  OAI22_X1 U459 ( .A1(n223), .A2(n194), .B1(n193), .B2(n303), .ZN(n159) );
  OAI22_X1 U460 ( .A1(n328), .A2(n196), .B1(n195), .B2(n303), .ZN(n161) );
  OAI22_X1 U461 ( .A1(n328), .A2(n231), .B1(n199), .B2(n303), .ZN(n139) );
  OAI22_X1 U462 ( .A1(n328), .A2(n197), .B1(n196), .B2(n304), .ZN(n162) );
  OAI22_X1 U463 ( .A1(n223), .A2(n192), .B1(n191), .B2(n303), .ZN(n99) );
  OAI22_X1 U464 ( .A1(n223), .A2(n191), .B1(n191), .B2(n304), .ZN(n131) );
  XNOR2_X1 U465 ( .A(n329), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U466 ( .A(n329), .B(b[6]), .ZN(n201) );
  INV_X1 U467 ( .A(n304), .ZN(n132) );
  OAI22_X1 U468 ( .A1(n328), .A2(n198), .B1(n197), .B2(n303), .ZN(n163) );
  XNOR2_X1 U469 ( .A(n329), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U470 ( .A(n329), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U471 ( .A(n330), .B(n329), .ZN(n207) );
  XNOR2_X1 U472 ( .A(n329), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U473 ( .A(n329), .B(b[3]), .ZN(n204) );
  INV_X1 U474 ( .A(n236), .ZN(n232) );
  XNOR2_X1 U475 ( .A(n329), .B(b[1]), .ZN(n206) );
  XOR2_X1 U476 ( .A(n236), .B(n135), .Z(n220) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70,
         n73, n74, n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n128, n129, n131, n132, n134, n135, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n229, n230, n231, n232, n233, n234, n235, n236,
         n244, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n289), .B(n150), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n100), .B(n151), .CI(n145), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n166), .B(n159), .CI(n153), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n170), .B(n163), .CO(n123), .S(n124) );
  OAI21_X1 U237 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  BUF_X1 U238 ( .A(n234), .Z(n327) );
  BUF_X1 U239 ( .A(n234), .Z(n280) );
  INV_X1 U240 ( .A(n290), .ZN(n287) );
  OR2_X1 U241 ( .A1(n172), .A2(n140), .ZN(n274) );
  XOR2_X1 U242 ( .A(n233), .B(a[6]), .Z(n275) );
  NOR2_X2 U243 ( .A1(n108), .A2(n113), .ZN(n44) );
  XOR2_X1 U244 ( .A(n168), .B(n161), .Z(n276) );
  XOR2_X1 U245 ( .A(n120), .B(n276), .Z(n118) );
  NAND2_X1 U246 ( .A1(n120), .A2(n168), .ZN(n277) );
  NAND2_X1 U247 ( .A1(n120), .A2(n161), .ZN(n278) );
  NAND2_X1 U248 ( .A1(n168), .A2(n161), .ZN(n279) );
  NAND3_X1 U249 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n117) );
  XOR2_X1 U250 ( .A(n290), .B(b[7]), .Z(n191) );
  INV_X1 U251 ( .A(n290), .ZN(n291) );
  CLKBUF_X1 U252 ( .A(n45), .Z(n281) );
  XNOR2_X1 U253 ( .A(n104), .B(n282), .ZN(n102) );
  XNOR2_X1 U254 ( .A(n109), .B(n106), .ZN(n282) );
  INV_X1 U255 ( .A(n34), .ZN(n283) );
  CLKBUF_X1 U256 ( .A(n216), .Z(n314) );
  CLKBUF_X1 U257 ( .A(n216), .Z(n334) );
  XOR2_X1 U258 ( .A(n236), .B(n135), .Z(n220) );
  AOI21_X1 U259 ( .B1(n321), .B2(n55), .A(n52), .ZN(n284) );
  AOI21_X1 U260 ( .B1(n321), .B2(n55), .A(n52), .ZN(n50) );
  XOR2_X1 U261 ( .A(n230), .B(b[6]), .Z(n183) );
  CLKBUF_X1 U262 ( .A(n296), .Z(n285) );
  XNOR2_X1 U263 ( .A(n158), .B(n146), .ZN(n106) );
  XOR2_X1 U264 ( .A(n327), .B(a[4]), .Z(n286) );
  OAI21_X1 U265 ( .B1(n285), .B2(n283), .A(n31), .ZN(n288) );
  OAI22_X1 U266 ( .A1(n223), .A2(n192), .B1(n191), .B2(n323), .ZN(n289) );
  INV_X1 U267 ( .A(n235), .ZN(n290) );
  CLKBUF_X3 U268 ( .A(n236), .Z(n322) );
  NOR2_X1 U269 ( .A1(n35), .A2(n30), .ZN(n292) );
  NAND2_X1 U270 ( .A1(n104), .A2(n109), .ZN(n293) );
  NAND2_X1 U271 ( .A1(n104), .A2(n106), .ZN(n294) );
  NAND2_X1 U272 ( .A1(n109), .A2(n106), .ZN(n295) );
  NAND3_X1 U273 ( .A1(n293), .A2(n294), .A3(n295), .ZN(n101) );
  NOR2_X1 U274 ( .A1(n92), .A2(n95), .ZN(n296) );
  CLKBUF_X1 U275 ( .A(n39), .Z(n297) );
  NOR2_X1 U276 ( .A1(n92), .A2(n95), .ZN(n30) );
  XNOR2_X1 U277 ( .A(n303), .B(n298), .ZN(product[14]) );
  XNOR2_X1 U278 ( .A(n141), .B(n83), .ZN(n298) );
  CLKBUF_X1 U279 ( .A(n330), .Z(n324) );
  NAND2_X2 U280 ( .A1(n220), .A2(n244), .ZN(n224) );
  BUF_X2 U281 ( .A(n330), .Z(n323) );
  CLKBUF_X1 U282 ( .A(n226), .Z(n325) );
  BUF_X1 U283 ( .A(n226), .Z(n326) );
  AND3_X1 U284 ( .A1(n309), .A2(n310), .A3(n308), .ZN(product[15]) );
  CLKBUF_X1 U285 ( .A(n70), .Z(n300) );
  NAND2_X1 U286 ( .A1(n219), .A2(n330), .ZN(n301) );
  NAND2_X1 U287 ( .A1(n219), .A2(n330), .ZN(n302) );
  NAND2_X1 U288 ( .A1(n330), .A2(n219), .ZN(n223) );
  NAND3_X1 U289 ( .A1(n307), .A2(n306), .A3(n305), .ZN(n303) );
  XOR2_X1 U290 ( .A(n85), .B(n84), .Z(n304) );
  XOR2_X1 U291 ( .A(n304), .B(n300), .Z(product[13]) );
  NAND2_X1 U292 ( .A1(n85), .A2(n84), .ZN(n305) );
  NAND2_X1 U293 ( .A1(n70), .A2(n85), .ZN(n306) );
  NAND2_X1 U294 ( .A1(n84), .A2(n70), .ZN(n307) );
  NAND3_X1 U295 ( .A1(n306), .A2(n305), .A3(n307), .ZN(n14) );
  NAND2_X1 U296 ( .A1(n141), .A2(n83), .ZN(n308) );
  NAND2_X1 U297 ( .A1(n303), .A2(n141), .ZN(n309) );
  NAND2_X1 U298 ( .A1(n83), .A2(n14), .ZN(n310) );
  CLKBUF_X1 U299 ( .A(n47), .Z(n311) );
  CLKBUF_X1 U300 ( .A(n20), .Z(n312) );
  NOR2_X1 U301 ( .A1(n102), .A2(n107), .ZN(n313) );
  AOI21_X1 U302 ( .B1(n297), .B2(n311), .A(n40), .ZN(n315) );
  NAND2_X1 U303 ( .A1(n217), .A2(n331), .ZN(n316) );
  XNOR2_X1 U304 ( .A(n234), .B(a[6]), .ZN(n225) );
  INV_X1 U305 ( .A(n35), .ZN(n74) );
  XNOR2_X1 U306 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U307 ( .A1(n74), .A2(n283), .ZN(n4) );
  INV_X1 U308 ( .A(n36), .ZN(n34) );
  INV_X1 U309 ( .A(n54), .ZN(n52) );
  INV_X1 U310 ( .A(n26), .ZN(n24) );
  AOI21_X1 U311 ( .B1(n318), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U312 ( .A(n66), .ZN(n64) );
  NAND2_X1 U313 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U314 ( .A(n48), .ZN(n77) );
  INV_X1 U315 ( .A(n69), .ZN(n67) );
  NOR2_X1 U316 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U317 ( .A1(n321), .A2(n54), .ZN(n8) );
  NAND2_X1 U318 ( .A1(n320), .A2(n19), .ZN(n1) );
  XOR2_X1 U319 ( .A(n10), .B(n62), .Z(product[3]) );
  NAND2_X1 U320 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U321 ( .A(n60), .ZN(n80) );
  XOR2_X1 U322 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U323 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U324 ( .A(n56), .ZN(n79) );
  XOR2_X1 U325 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U326 ( .A1(n31), .A2(n73), .ZN(n3) );
  AOI21_X1 U327 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U328 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U329 ( .A1(n76), .A2(n281), .ZN(n6) );
  INV_X1 U330 ( .A(n44), .ZN(n76) );
  XOR2_X1 U331 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U332 ( .A1(n319), .A2(n26), .ZN(n2) );
  NOR2_X1 U333 ( .A1(n35), .A2(n30), .ZN(n28) );
  NAND2_X1 U334 ( .A1(n96), .A2(n101), .ZN(n36) );
  XNOR2_X1 U335 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U336 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U337 ( .B1(n46), .B2(n44), .A(n281), .ZN(n43) );
  NAND2_X1 U338 ( .A1(n102), .A2(n107), .ZN(n42) );
  INV_X1 U339 ( .A(n59), .ZN(n58) );
  OAI21_X1 U340 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  XNOR2_X1 U341 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U342 ( .A1(n318), .A2(n66), .ZN(n11) );
  INV_X1 U343 ( .A(n19), .ZN(n17) );
  OR2_X1 U344 ( .A1(n158), .A2(n146), .ZN(n105) );
  AND2_X1 U345 ( .A1(n274), .A2(n69), .ZN(product[1]) );
  NOR2_X1 U346 ( .A1(n124), .A2(n139), .ZN(n60) );
  OR2_X1 U347 ( .A1(n171), .A2(n164), .ZN(n318) );
  NAND2_X1 U348 ( .A1(n108), .A2(n113), .ZN(n45) );
  NOR2_X1 U349 ( .A1(n122), .A2(n123), .ZN(n56) );
  NOR2_X1 U350 ( .A1(n114), .A2(n117), .ZN(n48) );
  INV_X1 U351 ( .A(n83), .ZN(n84) );
  OR2_X1 U352 ( .A1(n88), .A2(n91), .ZN(n319) );
  NAND2_X1 U353 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U354 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U355 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U356 ( .A1(n122), .A2(n123), .ZN(n57) );
  NAND2_X1 U357 ( .A1(n92), .A2(n95), .ZN(n31) );
  OR2_X1 U358 ( .A1(n87), .A2(n86), .ZN(n320) );
  OR2_X1 U359 ( .A1(n118), .A2(n121), .ZN(n321) );
  OR2_X1 U360 ( .A1(n314), .A2(n231), .ZN(n199) );
  OAI22_X1 U361 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  AND2_X1 U362 ( .A1(n314), .A2(n126), .ZN(n148) );
  OR2_X1 U363 ( .A1(n334), .A2(n229), .ZN(n181) );
  OR2_X1 U364 ( .A1(n334), .A2(n230), .ZN(n190) );
  INV_X1 U365 ( .A(n128), .ZN(n149) );
  INV_X1 U366 ( .A(n89), .ZN(n90) );
  AND2_X1 U367 ( .A1(n334), .A2(n129), .ZN(n156) );
  OAI22_X1 U368 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U369 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  OR2_X1 U370 ( .A1(n314), .A2(n232), .ZN(n208) );
  OAI22_X1 U371 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U372 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  BUF_X1 U373 ( .A(n225), .Z(n333) );
  INV_X1 U374 ( .A(n125), .ZN(n141) );
  AND2_X1 U375 ( .A1(n334), .A2(n132), .ZN(n164) );
  NAND2_X1 U376 ( .A1(n275), .A2(n331), .ZN(n221) );
  AND2_X1 U377 ( .A1(n216), .A2(n135), .ZN(product[0]) );
  XNOR2_X1 U378 ( .A(n235), .B(a[4]), .ZN(n226) );
  BUF_X1 U379 ( .A(n225), .Z(n332) );
  OAI22_X1 U380 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U381 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  NAND2_X1 U382 ( .A1(n171), .A2(n164), .ZN(n66) );
  OAI22_X1 U383 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  NAND2_X1 U384 ( .A1(n286), .A2(n326), .ZN(n328) );
  NAND2_X1 U385 ( .A1(n218), .A2(n226), .ZN(n329) );
  NAND2_X1 U386 ( .A1(n286), .A2(n226), .ZN(n222) );
  XNOR2_X1 U387 ( .A(n236), .B(a[2]), .ZN(n330) );
  INV_X1 U388 ( .A(n134), .ZN(n165) );
  XNOR2_X1 U389 ( .A(n314), .B(n233), .ZN(n180) );
  XNOR2_X1 U390 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U391 ( .A(n233), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U392 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U393 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U394 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U395 ( .A(b[7]), .B(n233), .ZN(n173) );
  INV_X1 U396 ( .A(n233), .ZN(n229) );
  XOR2_X1 U397 ( .A(n233), .B(a[6]), .Z(n217) );
  INV_X1 U398 ( .A(n99), .ZN(n100) );
  AOI21_X1 U399 ( .B1(n37), .B2(n292), .A(n288), .ZN(n27) );
  INV_X1 U400 ( .A(n291), .ZN(n231) );
  XNOR2_X1 U401 ( .A(n291), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U402 ( .A(n287), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U403 ( .A(n291), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U404 ( .A(n287), .B(b[5]), .ZN(n193) );
  INV_X1 U405 ( .A(n131), .ZN(n157) );
  NAND2_X1 U406 ( .A1(n124), .A2(n139), .ZN(n61) );
  BUF_X1 U407 ( .A(n225), .Z(n331) );
  NAND2_X1 U408 ( .A1(n118), .A2(n121), .ZN(n54) );
  NOR2_X1 U409 ( .A1(n102), .A2(n107), .ZN(n41) );
  OAI22_X1 U410 ( .A1(n224), .A2(n200), .B1(n200), .B2(n244), .ZN(n134) );
  XOR2_X1 U411 ( .A(n235), .B(a[2]), .Z(n219) );
  XNOR2_X1 U412 ( .A(n334), .B(n287), .ZN(n198) );
  XNOR2_X1 U413 ( .A(n287), .B(b[6]), .ZN(n192) );
  OAI21_X1 U414 ( .B1(n296), .B2(n36), .A(n31), .ZN(n29) );
  INV_X1 U415 ( .A(n30), .ZN(n73) );
  OAI21_X1 U416 ( .B1(n48), .B2(n50), .A(n49), .ZN(n47) );
  AOI21_X1 U417 ( .B1(n29), .B2(n319), .A(n24), .ZN(n22) );
  NAND2_X1 U418 ( .A1(n28), .A2(n319), .ZN(n21) );
  INV_X1 U419 ( .A(n313), .ZN(n75) );
  OAI22_X1 U420 ( .A1(n173), .A2(n316), .B1(n173), .B2(n332), .ZN(n125) );
  OAI21_X1 U421 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  OAI22_X1 U422 ( .A1(n316), .A2(n174), .B1(n173), .B2(n333), .ZN(n83) );
  NOR2_X1 U423 ( .A1(n313), .A2(n44), .ZN(n39) );
  OAI21_X1 U424 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI22_X1 U425 ( .A1(n316), .A2(n175), .B1(n174), .B2(n332), .ZN(n142) );
  OAI22_X1 U426 ( .A1(n316), .A2(n176), .B1(n175), .B2(n333), .ZN(n143) );
  OAI22_X1 U427 ( .A1(n316), .A2(n177), .B1(n176), .B2(n332), .ZN(n144) );
  INV_X1 U428 ( .A(n333), .ZN(n126) );
  OAI22_X1 U429 ( .A1(n316), .A2(n178), .B1(n177), .B2(n332), .ZN(n145) );
  OAI22_X1 U430 ( .A1(n316), .A2(n179), .B1(n178), .B2(n333), .ZN(n146) );
  OAI22_X1 U431 ( .A1(n221), .A2(n229), .B1(n181), .B2(n332), .ZN(n137) );
  OAI22_X1 U432 ( .A1(n221), .A2(n180), .B1(n179), .B2(n333), .ZN(n147) );
  XNOR2_X1 U433 ( .A(n55), .B(n8), .ZN(product[5]) );
  INV_X1 U434 ( .A(n311), .ZN(n46) );
  AOI21_X1 U435 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U436 ( .A1(n140), .A2(n172), .ZN(n69) );
  XNOR2_X1 U437 ( .A(n322), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U438 ( .A(n322), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U439 ( .A(n322), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U440 ( .A(n322), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U441 ( .A(n322), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U442 ( .A(n322), .B(b[3]), .ZN(n204) );
  XNOR2_X1 U443 ( .A(n314), .B(n322), .ZN(n207) );
  INV_X1 U444 ( .A(n322), .ZN(n232) );
  XOR2_X1 U445 ( .A(n7), .B(n284), .Z(product[6]) );
  OAI22_X1 U446 ( .A1(n182), .A2(n328), .B1(n182), .B2(n325), .ZN(n128) );
  OAI22_X1 U447 ( .A1(n328), .A2(n188), .B1(n187), .B2(n326), .ZN(n154) );
  OAI22_X1 U448 ( .A1(n328), .A2(n183), .B1(n182), .B2(n325), .ZN(n89) );
  OAI22_X1 U449 ( .A1(n329), .A2(n185), .B1(n184), .B2(n326), .ZN(n151) );
  OAI22_X1 U450 ( .A1(n329), .A2(n187), .B1(n186), .B2(n325), .ZN(n153) );
  OAI22_X1 U451 ( .A1(n329), .A2(n184), .B1(n183), .B2(n326), .ZN(n150) );
  OAI22_X1 U452 ( .A1(n329), .A2(n186), .B1(n185), .B2(n326), .ZN(n152) );
  INV_X1 U453 ( .A(n326), .ZN(n129) );
  OAI22_X1 U454 ( .A1(n222), .A2(n230), .B1(n190), .B2(n325), .ZN(n138) );
  OAI22_X1 U455 ( .A1(n222), .A2(n189), .B1(n188), .B2(n325), .ZN(n155) );
  INV_X1 U456 ( .A(n15), .ZN(n70) );
  XNOR2_X1 U457 ( .A(n280), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U458 ( .A(n280), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U459 ( .A(n280), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U460 ( .A(n280), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U461 ( .A(n280), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U462 ( .A(n334), .B(n280), .ZN(n189) );
  INV_X1 U463 ( .A(n327), .ZN(n230) );
  XOR2_X1 U464 ( .A(n327), .B(a[4]), .Z(n218) );
  XNOR2_X1 U465 ( .A(n233), .B(b[1]), .ZN(n179) );
  XNOR2_X1 U466 ( .A(n280), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U467 ( .A(n291), .B(b[1]), .ZN(n197) );
  XNOR2_X1 U468 ( .A(n322), .B(b[1]), .ZN(n206) );
  XNOR2_X1 U469 ( .A(n312), .B(n1), .ZN(product[12]) );
  INV_X1 U470 ( .A(n315), .ZN(n37) );
  AOI21_X1 U471 ( .B1(n20), .B2(n320), .A(n17), .ZN(n15) );
  OAI22_X1 U472 ( .A1(n302), .A2(n193), .B1(n192), .B2(n324), .ZN(n158) );
  OAI22_X1 U473 ( .A1(n301), .A2(n195), .B1(n194), .B2(n323), .ZN(n160) );
  OAI22_X1 U474 ( .A1(n302), .A2(n194), .B1(n193), .B2(n324), .ZN(n159) );
  OAI22_X1 U475 ( .A1(n301), .A2(n196), .B1(n195), .B2(n324), .ZN(n161) );
  OAI22_X1 U476 ( .A1(n301), .A2(n231), .B1(n199), .B2(n323), .ZN(n139) );
  OAI22_X1 U477 ( .A1(n302), .A2(n197), .B1(n196), .B2(n323), .ZN(n162) );
  OAI22_X1 U478 ( .A1(n223), .A2(n192), .B1(n191), .B2(n323), .ZN(n99) );
  OAI22_X1 U479 ( .A1(n191), .A2(n223), .B1(n191), .B2(n323), .ZN(n131) );
  INV_X1 U480 ( .A(n323), .ZN(n132) );
  OAI22_X1 U481 ( .A1(n301), .A2(n198), .B1(n197), .B2(n324), .ZN(n163) );
  INV_X2 U482 ( .A(n135), .ZN(n244) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n73,
         n74, n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n128, n129, n131, n132, n134, n135, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n229, n230, n231, n232, n233, n234, n235, n236,
         n244, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n150), .B(n283), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n145), .B(n100), .CI(n151), .CO(n97), .S(n98) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n159), .B(n166), .CI(n153), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n167), .B(n148), .CI(n160), .CO(n115), .S(n116) );
  HA_X1 U115 ( .A(n155), .B(n138), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  BUF_X2 U237 ( .A(n216), .Z(n337) );
  OR2_X1 U238 ( .A1(n172), .A2(n140), .ZN(n274) );
  XNOR2_X1 U239 ( .A(n280), .B(b[7]), .ZN(n275) );
  AND2_X1 U240 ( .A1(n96), .A2(n101), .ZN(n276) );
  CLKBUF_X1 U241 ( .A(b[4]), .Z(n277) );
  NOR2_X2 U242 ( .A1(n114), .A2(n117), .ZN(n48) );
  CLKBUF_X1 U243 ( .A(n28), .Z(n278) );
  CLKBUF_X1 U244 ( .A(n236), .Z(n279) );
  CLKBUF_X3 U245 ( .A(n235), .Z(n280) );
  CLKBUF_X1 U246 ( .A(n236), .Z(n281) );
  NAND3_X1 U247 ( .A1(n303), .A2(n304), .A3(n305), .ZN(n282) );
  OAI22_X1 U248 ( .A1(n297), .A2(n192), .B1(n191), .B2(n336), .ZN(n283) );
  NOR2_X1 U249 ( .A1(n92), .A2(n95), .ZN(n284) );
  NOR2_X1 U250 ( .A1(n92), .A2(n95), .ZN(n30) );
  AND3_X1 U251 ( .A1(n307), .A2(n308), .A3(n309), .ZN(product[15]) );
  XOR2_X1 U252 ( .A(n161), .B(n168), .Z(n286) );
  XOR2_X1 U253 ( .A(n120), .B(n286), .Z(n118) );
  NAND2_X1 U254 ( .A1(n120), .A2(n161), .ZN(n287) );
  NAND2_X1 U255 ( .A1(n120), .A2(n168), .ZN(n288) );
  NAND2_X1 U256 ( .A1(n161), .A2(n168), .ZN(n289) );
  NAND3_X1 U257 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n117) );
  NAND2_X1 U258 ( .A1(n220), .A2(n244), .ZN(n290) );
  NAND2_X1 U259 ( .A1(n220), .A2(n244), .ZN(n291) );
  NAND2_X1 U260 ( .A1(n220), .A2(n244), .ZN(n224) );
  INV_X1 U261 ( .A(n276), .ZN(n292) );
  CLKBUF_X1 U262 ( .A(n221), .Z(n322) );
  NAND2_X1 U263 ( .A1(n236), .A2(n294), .ZN(n295) );
  NAND2_X1 U264 ( .A1(n293), .A2(n135), .ZN(n296) );
  NAND2_X1 U265 ( .A1(n295), .A2(n296), .ZN(n220) );
  INV_X1 U266 ( .A(n236), .ZN(n293) );
  INV_X1 U267 ( .A(n135), .ZN(n294) );
  NAND2_X1 U268 ( .A1(n227), .A2(n219), .ZN(n297) );
  NAND2_X1 U269 ( .A1(n227), .A2(n219), .ZN(n223) );
  NAND2_X1 U270 ( .A1(n218), .A2(n226), .ZN(n298) );
  NAND2_X1 U271 ( .A1(n218), .A2(n226), .ZN(n299) );
  NAND2_X1 U272 ( .A1(n218), .A2(n226), .ZN(n222) );
  CLKBUF_X1 U273 ( .A(n70), .Z(n300) );
  XNOR2_X1 U274 ( .A(n301), .B(n111), .ZN(n104) );
  XNOR2_X1 U275 ( .A(n165), .B(n152), .ZN(n301) );
  XOR2_X1 U276 ( .A(n85), .B(n84), .Z(n302) );
  XOR2_X1 U277 ( .A(n302), .B(n300), .Z(product[13]) );
  NAND2_X1 U278 ( .A1(n85), .A2(n84), .ZN(n303) );
  NAND2_X1 U279 ( .A1(n70), .A2(n85), .ZN(n304) );
  NAND2_X1 U280 ( .A1(n70), .A2(n84), .ZN(n305) );
  NAND3_X1 U281 ( .A1(n303), .A2(n304), .A3(n305), .ZN(n14) );
  XOR2_X1 U282 ( .A(n141), .B(n83), .Z(n306) );
  XOR2_X1 U283 ( .A(n306), .B(n282), .Z(product[14]) );
  NAND2_X1 U284 ( .A1(n141), .A2(n83), .ZN(n307) );
  NAND2_X1 U285 ( .A1(n14), .A2(n141), .ZN(n308) );
  NAND2_X1 U286 ( .A1(n14), .A2(n83), .ZN(n309) );
  XOR2_X1 U287 ( .A(n109), .B(n106), .Z(n310) );
  XOR2_X1 U288 ( .A(n310), .B(n104), .Z(n102) );
  NAND2_X1 U289 ( .A1(n165), .A2(n152), .ZN(n311) );
  NAND2_X1 U290 ( .A1(n165), .A2(n111), .ZN(n312) );
  NAND2_X1 U291 ( .A1(n152), .A2(n111), .ZN(n313) );
  NAND3_X1 U292 ( .A1(n311), .A2(n312), .A3(n313), .ZN(n103) );
  NAND2_X1 U293 ( .A1(n109), .A2(n106), .ZN(n314) );
  NAND2_X1 U294 ( .A1(n109), .A2(n104), .ZN(n315) );
  NAND2_X1 U295 ( .A1(n106), .A2(n104), .ZN(n316) );
  NAND3_X1 U296 ( .A1(n314), .A2(n315), .A3(n316), .ZN(n101) );
  AOI21_X1 U297 ( .B1(n327), .B2(n55), .A(n52), .ZN(n317) );
  AOI21_X1 U298 ( .B1(n327), .B2(n55), .A(n52), .ZN(n50) );
  BUF_X2 U299 ( .A(n226), .Z(n328) );
  CLKBUF_X1 U300 ( .A(n20), .Z(n318) );
  CLKBUF_X1 U301 ( .A(n234), .Z(n319) );
  OAI21_X1 U302 ( .B1(n48), .B2(n317), .A(n49), .ZN(n320) );
  AOI21_X1 U303 ( .B1(n39), .B2(n320), .A(n40), .ZN(n321) );
  INV_X1 U304 ( .A(n35), .ZN(n74) );
  INV_X1 U305 ( .A(n320), .ZN(n46) );
  XNOR2_X1 U306 ( .A(n37), .B(n4), .ZN(product[9]) );
  NAND2_X1 U307 ( .A1(n74), .A2(n292), .ZN(n4) );
  INV_X1 U308 ( .A(n66), .ZN(n64) );
  INV_X1 U309 ( .A(n26), .ZN(n24) );
  OAI21_X1 U310 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  INV_X1 U311 ( .A(n59), .ZN(n58) );
  NOR2_X1 U312 ( .A1(n96), .A2(n101), .ZN(n35) );
  NAND2_X1 U313 ( .A1(n325), .A2(n19), .ZN(n1) );
  XOR2_X1 U314 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U315 ( .A1(n76), .A2(n45), .ZN(n6) );
  INV_X1 U316 ( .A(n44), .ZN(n76) );
  XOR2_X1 U317 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U318 ( .A1(n73), .A2(n31), .ZN(n3) );
  AOI21_X1 U319 ( .B1(n37), .B2(n74), .A(n276), .ZN(n32) );
  XOR2_X1 U320 ( .A(n27), .B(n2), .Z(product[11]) );
  NAND2_X1 U321 ( .A1(n323), .A2(n26), .ZN(n2) );
  XNOR2_X1 U322 ( .A(n8), .B(n55), .ZN(product[5]) );
  XNOR2_X1 U323 ( .A(n43), .B(n5), .ZN(product[8]) );
  OAI21_X1 U324 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U325 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U326 ( .A1(n324), .A2(n66), .ZN(n11) );
  INV_X1 U327 ( .A(n69), .ZN(n67) );
  XOR2_X1 U328 ( .A(n10), .B(n62), .Z(product[3]) );
  NAND2_X1 U329 ( .A1(n80), .A2(n61), .ZN(n10) );
  INV_X1 U330 ( .A(n60), .ZN(n80) );
  NAND2_X1 U331 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U332 ( .A(n48), .ZN(n77) );
  XOR2_X1 U333 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U334 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U335 ( .A(n56), .ZN(n79) );
  INV_X1 U336 ( .A(n19), .ZN(n17) );
  NOR2_X1 U337 ( .A1(n108), .A2(n113), .ZN(n44) );
  XNOR2_X1 U338 ( .A(n158), .B(n146), .ZN(n106) );
  OR2_X1 U339 ( .A1(n158), .A2(n146), .ZN(n105) );
  NOR2_X1 U340 ( .A1(n122), .A2(n123), .ZN(n56) );
  INV_X1 U341 ( .A(n83), .ZN(n84) );
  OR2_X1 U342 ( .A1(n88), .A2(n91), .ZN(n323) );
  NAND2_X1 U343 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U344 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U345 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U346 ( .A1(n122), .A2(n123), .ZN(n57) );
  OR2_X1 U347 ( .A1(n171), .A2(n164), .ZN(n324) );
  OR2_X1 U348 ( .A1(n87), .A2(n86), .ZN(n325) );
  AND2_X1 U349 ( .A1(n274), .A2(n69), .ZN(product[1]) );
  OR2_X1 U350 ( .A1(n118), .A2(n121), .ZN(n327) );
  OR2_X1 U351 ( .A1(n337), .A2(n231), .ZN(n199) );
  OR2_X1 U352 ( .A1(n337), .A2(n232), .ZN(n208) );
  INV_X1 U353 ( .A(n128), .ZN(n149) );
  INV_X1 U354 ( .A(n89), .ZN(n90) );
  AND2_X1 U355 ( .A1(n337), .A2(n129), .ZN(n156) );
  OAI22_X1 U356 ( .A1(n291), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OR2_X1 U357 ( .A1(n337), .A2(n230), .ZN(n190) );
  AND2_X1 U358 ( .A1(n337), .A2(n126), .ZN(n148) );
  BUF_X1 U359 ( .A(n225), .Z(n331) );
  BUF_X1 U360 ( .A(n225), .Z(n330) );
  INV_X1 U361 ( .A(n125), .ZN(n141) );
  INV_X1 U362 ( .A(n131), .ZN(n157) );
  AND2_X1 U363 ( .A1(n337), .A2(n132), .ZN(n164) );
  OR2_X1 U364 ( .A1(n337), .A2(n229), .ZN(n181) );
  INV_X1 U365 ( .A(n135), .ZN(n244) );
  NAND2_X1 U366 ( .A1(n217), .A2(n329), .ZN(n221) );
  AND2_X1 U367 ( .A1(n337), .A2(n135), .ZN(product[0]) );
  NAND2_X1 U368 ( .A1(n171), .A2(n164), .ZN(n66) );
  OAI22_X1 U369 ( .A1(n290), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  XNOR2_X1 U370 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U371 ( .A(n233), .B(n277), .ZN(n176) );
  XNOR2_X1 U372 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U373 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U374 ( .A(n337), .B(n233), .ZN(n180) );
  INV_X1 U375 ( .A(n233), .ZN(n229) );
  XNOR2_X1 U376 ( .A(n235), .B(a[4]), .ZN(n226) );
  BUF_X1 U377 ( .A(n225), .Z(n329) );
  XNOR2_X1 U378 ( .A(n234), .B(a[6]), .ZN(n225) );
  OAI22_X1 U379 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OAI22_X1 U380 ( .A1(n290), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  NAND2_X1 U381 ( .A1(n75), .A2(n42), .ZN(n5) );
  INV_X1 U382 ( .A(n134), .ZN(n165) );
  NAND2_X1 U383 ( .A1(n108), .A2(n113), .ZN(n45) );
  NAND2_X1 U384 ( .A1(n102), .A2(n107), .ZN(n42) );
  XOR2_X1 U385 ( .A(n233), .B(a[6]), .Z(n217) );
  NOR2_X1 U386 ( .A1(n102), .A2(n107), .ZN(n332) );
  NOR2_X1 U387 ( .A1(n102), .A2(n107), .ZN(n41) );
  CLKBUF_X1 U388 ( .A(n234), .Z(n333) );
  NAND2_X1 U389 ( .A1(n327), .A2(n54), .ZN(n8) );
  INV_X1 U390 ( .A(n54), .ZN(n52) );
  CLKBUF_X1 U391 ( .A(n29), .Z(n334) );
  XNOR2_X1 U392 ( .A(n236), .B(a[2]), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n236), .B(a[2]), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n236), .B(a[2]), .ZN(n227) );
  NAND2_X1 U395 ( .A1(n28), .A2(n323), .ZN(n21) );
  OAI21_X1 U396 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  NOR2_X1 U397 ( .A1(n35), .A2(n284), .ZN(n28) );
  NAND2_X1 U398 ( .A1(n96), .A2(n101), .ZN(n36) );
  XNOR2_X1 U399 ( .A(n333), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U400 ( .A(n319), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U401 ( .A(n319), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U402 ( .A(n337), .B(n319), .ZN(n189) );
  XNOR2_X1 U403 ( .A(n333), .B(b[5]), .ZN(n184) );
  INV_X1 U404 ( .A(n234), .ZN(n230) );
  XOR2_X1 U405 ( .A(n234), .B(a[4]), .Z(n218) );
  NAND2_X1 U406 ( .A1(n124), .A2(n139), .ZN(n61) );
  NOR2_X1 U407 ( .A1(n124), .A2(n139), .ZN(n60) );
  OAI22_X1 U408 ( .A1(n291), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U409 ( .A1(n291), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  XNOR2_X1 U410 ( .A(n319), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U411 ( .A(n233), .B(b[3]), .ZN(n177) );
  XOR2_X1 U412 ( .A(n7), .B(n317), .Z(product[6]) );
  INV_X1 U413 ( .A(n99), .ZN(n100) );
  AOI21_X1 U414 ( .B1(n29), .B2(n323), .A(n24), .ZN(n22) );
  AOI21_X1 U415 ( .B1(n37), .B2(n278), .A(n334), .ZN(n27) );
  NAND2_X1 U416 ( .A1(n172), .A2(n140), .ZN(n69) );
  AOI21_X1 U417 ( .B1(n324), .B2(n67), .A(n64), .ZN(n62) );
  OAI21_X1 U418 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  OAI22_X1 U419 ( .A1(n290), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  XNOR2_X1 U420 ( .A(n319), .B(b[1]), .ZN(n188) );
  XNOR2_X1 U421 ( .A(n233), .B(b[1]), .ZN(n179) );
  INV_X1 U422 ( .A(n332), .ZN(n75) );
  NOR2_X1 U423 ( .A1(n332), .A2(n44), .ZN(n39) );
  OAI21_X1 U424 ( .B1(n45), .B2(n41), .A(n42), .ZN(n40) );
  XNOR2_X1 U425 ( .A(n233), .B(b[7]), .ZN(n173) );
  XNOR2_X1 U426 ( .A(n333), .B(b[7]), .ZN(n182) );
  OAI22_X1 U427 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U428 ( .A1(n200), .A2(n290), .B1(n200), .B2(n244), .ZN(n134) );
  NAND2_X1 U429 ( .A1(n118), .A2(n121), .ZN(n54) );
  OAI22_X1 U430 ( .A1(n182), .A2(n299), .B1(n182), .B2(n328), .ZN(n128) );
  OAI22_X1 U431 ( .A1(n222), .A2(n188), .B1(n187), .B2(n328), .ZN(n154) );
  OAI22_X1 U432 ( .A1(n298), .A2(n183), .B1(n182), .B2(n328), .ZN(n89) );
  OAI22_X1 U433 ( .A1(n298), .A2(n184), .B1(n183), .B2(n328), .ZN(n150) );
  INV_X1 U434 ( .A(n328), .ZN(n129) );
  OAI22_X1 U435 ( .A1(n222), .A2(n185), .B1(n184), .B2(n328), .ZN(n151) );
  OAI22_X1 U436 ( .A1(n299), .A2(n187), .B1(n186), .B2(n328), .ZN(n153) );
  OAI22_X1 U437 ( .A1(n222), .A2(n186), .B1(n185), .B2(n328), .ZN(n152) );
  OAI22_X1 U438 ( .A1(n222), .A2(n230), .B1(n190), .B2(n328), .ZN(n138) );
  OAI22_X1 U439 ( .A1(n299), .A2(n189), .B1(n188), .B2(n328), .ZN(n155) );
  XNOR2_X1 U440 ( .A(n280), .B(b[3]), .ZN(n195) );
  XNOR2_X1 U441 ( .A(n280), .B(b[2]), .ZN(n196) );
  XNOR2_X1 U442 ( .A(n280), .B(b[4]), .ZN(n194) );
  INV_X1 U443 ( .A(n280), .ZN(n231) );
  XNOR2_X1 U444 ( .A(n280), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U445 ( .A(n280), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U446 ( .A(n337), .B(n280), .ZN(n198) );
  XNOR2_X1 U447 ( .A(n280), .B(b[1]), .ZN(n197) );
  XOR2_X1 U448 ( .A(n235), .B(a[2]), .Z(n219) );
  INV_X1 U449 ( .A(n284), .ZN(n73) );
  NAND2_X1 U450 ( .A1(n92), .A2(n95), .ZN(n31) );
  INV_X1 U451 ( .A(n15), .ZN(n70) );
  XNOR2_X1 U452 ( .A(n280), .B(b[7]), .ZN(n191) );
  OAI22_X1 U453 ( .A1(n173), .A2(n322), .B1(n173), .B2(n330), .ZN(n125) );
  OAI22_X1 U454 ( .A1(n322), .A2(n174), .B1(n173), .B2(n331), .ZN(n83) );
  OAI22_X1 U455 ( .A1(n322), .A2(n175), .B1(n174), .B2(n330), .ZN(n142) );
  OAI22_X1 U456 ( .A1(n322), .A2(n176), .B1(n175), .B2(n330), .ZN(n143) );
  OAI22_X1 U457 ( .A1(n322), .A2(n177), .B1(n176), .B2(n331), .ZN(n144) );
  INV_X1 U458 ( .A(n331), .ZN(n126) );
  OAI22_X1 U459 ( .A1(n221), .A2(n179), .B1(n178), .B2(n331), .ZN(n146) );
  OAI22_X1 U460 ( .A1(n221), .A2(n178), .B1(n177), .B2(n330), .ZN(n145) );
  OAI22_X1 U461 ( .A1(n221), .A2(n229), .B1(n181), .B2(n330), .ZN(n137) );
  OAI22_X1 U462 ( .A1(n221), .A2(n180), .B1(n179), .B2(n331), .ZN(n147) );
  OAI21_X1 U463 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  OAI21_X1 U464 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U465 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  XNOR2_X1 U466 ( .A(n318), .B(n1), .ZN(product[12]) );
  INV_X1 U467 ( .A(n321), .ZN(n37) );
  AOI21_X1 U468 ( .B1(n20), .B2(n325), .A(n17), .ZN(n15) );
  OAI22_X1 U469 ( .A1(n223), .A2(n193), .B1(n192), .B2(n335), .ZN(n158) );
  OAI22_X1 U470 ( .A1(n223), .A2(n195), .B1(n194), .B2(n335), .ZN(n160) );
  OAI22_X1 U471 ( .A1(n297), .A2(n194), .B1(n193), .B2(n336), .ZN(n159) );
  OAI22_X1 U472 ( .A1(n223), .A2(n196), .B1(n195), .B2(n336), .ZN(n161) );
  OAI22_X1 U473 ( .A1(n223), .A2(n231), .B1(n199), .B2(n335), .ZN(n139) );
  OAI22_X1 U474 ( .A1(n223), .A2(n197), .B1(n196), .B2(n336), .ZN(n162) );
  OAI22_X1 U475 ( .A1(n297), .A2(n192), .B1(n191), .B2(n336), .ZN(n99) );
  OAI22_X1 U476 ( .A1(n275), .A2(n297), .B1(n275), .B2(n335), .ZN(n131) );
  XNOR2_X1 U477 ( .A(n279), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U478 ( .A(n236), .B(b[6]), .ZN(n201) );
  INV_X1 U479 ( .A(n336), .ZN(n132) );
  OAI22_X1 U480 ( .A1(n223), .A2(n198), .B1(n197), .B2(n335), .ZN(n163) );
  XNOR2_X1 U481 ( .A(n281), .B(n277), .ZN(n203) );
  XNOR2_X1 U482 ( .A(n236), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U483 ( .A(n337), .B(n281), .ZN(n207) );
  XNOR2_X1 U484 ( .A(n281), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U485 ( .A(n279), .B(b[3]), .ZN(n204) );
  INV_X1 U486 ( .A(n236), .ZN(n232) );
  XNOR2_X1 U487 ( .A(n281), .B(b[1]), .ZN(n206) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n14, n15, n17, n19, n20, n21,
         n22, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n64, n66, n67, n69, n70, n73,
         n74, n75, n76, n77, n79, n80, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n128, n129, n131, n132, n134, n135, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n216, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n229, n230, n231, n232, n233, n234, n235, n236, n244,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344;
  assign n135 = a[0];
  assign n216 = b[0];
  assign n233 = a[7];
  assign n234 = a[5];
  assign n235 = a[3];
  assign n236 = a[1];

  FA_X1 U97 ( .A(n142), .B(n89), .CI(n149), .CO(n85), .S(n86) );
  FA_X1 U98 ( .A(n90), .B(n143), .CI(n93), .CO(n87), .S(n88) );
  FA_X1 U100 ( .A(n97), .B(n144), .CI(n94), .CO(n91), .S(n92) );
  FA_X1 U101 ( .A(n150), .B(n322), .CI(n157), .CO(n93), .S(n94) );
  FA_X1 U102 ( .A(n103), .B(n105), .CI(n98), .CO(n95), .S(n96) );
  FA_X1 U103 ( .A(n100), .B(n151), .CI(n145), .CO(n97), .S(n98) );
  FA_X1 U106 ( .A(n165), .B(n152), .CI(n111), .CO(n103), .S(n104) );
  FA_X1 U109 ( .A(n115), .B(n112), .CI(n110), .CO(n107), .S(n108) );
  FA_X1 U110 ( .A(n159), .B(n153), .CI(n166), .CO(n109), .S(n110) );
  HA_X1 U111 ( .A(n147), .B(n137), .CO(n111), .S(n112) );
  FA_X1 U112 ( .A(n119), .B(n154), .CI(n116), .CO(n113), .S(n114) );
  FA_X1 U113 ( .A(n160), .B(n148), .CI(n167), .CO(n115), .S(n116) );
  HA_X1 U115 ( .A(n138), .B(n155), .CO(n119), .S(n120) );
  FA_X1 U116 ( .A(n169), .B(n156), .CI(n162), .CO(n121), .S(n122) );
  HA_X1 U117 ( .A(n163), .B(n170), .CO(n123), .S(n124) );
  OR2_X1 U237 ( .A1(n118), .A2(n121), .ZN(n333) );
  BUF_X2 U238 ( .A(n234), .Z(n335) );
  BUF_X2 U239 ( .A(n234), .Z(n293) );
  OAI22_X1 U240 ( .A1(n222), .A2(n189), .B1(n188), .B2(n338), .ZN(n155) );
  BUF_X2 U241 ( .A(n225), .Z(n336) );
  OR2_X1 U242 ( .A1(n172), .A2(n140), .ZN(n274) );
  XOR2_X1 U243 ( .A(n168), .B(n161), .Z(n275) );
  XOR2_X1 U244 ( .A(n120), .B(n275), .Z(n118) );
  NAND2_X1 U245 ( .A1(n120), .A2(n168), .ZN(n276) );
  NAND2_X1 U246 ( .A1(n120), .A2(n161), .ZN(n277) );
  NAND2_X1 U247 ( .A1(n168), .A2(n161), .ZN(n278) );
  NAND3_X1 U248 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n117) );
  CLKBUF_X1 U249 ( .A(n35), .Z(n279) );
  CLKBUF_X1 U250 ( .A(n235), .Z(n280) );
  XOR2_X1 U251 ( .A(n233), .B(a[6]), .Z(n281) );
  NAND2_X1 U252 ( .A1(n236), .A2(n283), .ZN(n284) );
  NAND2_X1 U253 ( .A1(n282), .A2(n135), .ZN(n285) );
  NAND2_X1 U254 ( .A1(n284), .A2(n285), .ZN(n220) );
  INV_X1 U255 ( .A(n236), .ZN(n282) );
  INV_X1 U256 ( .A(n135), .ZN(n283) );
  XNOR2_X1 U257 ( .A(n305), .B(n286), .ZN(product[14]) );
  XNOR2_X1 U258 ( .A(n141), .B(n83), .ZN(n286) );
  XOR2_X1 U259 ( .A(n335), .B(a[4]), .Z(n287) );
  XNOR2_X1 U260 ( .A(n235), .B(a[2]), .ZN(n288) );
  INV_X1 U261 ( .A(n288), .ZN(n313) );
  XNOR2_X1 U262 ( .A(n234), .B(a[6]), .ZN(n225) );
  AND2_X1 U263 ( .A1(n118), .A2(n121), .ZN(n52) );
  NAND2_X1 U264 ( .A1(n218), .A2(n226), .ZN(n289) );
  CLKBUF_X1 U265 ( .A(n236), .Z(n290) );
  INV_X1 U266 ( .A(n77), .ZN(n291) );
  NOR2_X1 U267 ( .A1(n114), .A2(n117), .ZN(n48) );
  CLKBUF_X1 U268 ( .A(n44), .Z(n292) );
  BUF_X1 U269 ( .A(n225), .Z(n294) );
  XNOR2_X1 U270 ( .A(n104), .B(n295), .ZN(n102) );
  XNOR2_X1 U271 ( .A(n109), .B(n106), .ZN(n295) );
  BUF_X2 U272 ( .A(n317), .Z(n296) );
  CLKBUF_X1 U273 ( .A(n235), .Z(n297) );
  CLKBUF_X1 U274 ( .A(n289), .Z(n298) );
  AND3_X1 U275 ( .A1(n311), .A2(n312), .A3(n310), .ZN(product[15]) );
  CLKBUF_X1 U276 ( .A(n45), .Z(n300) );
  XNOR2_X1 U277 ( .A(n235), .B(a[4]), .ZN(n301) );
  CLKBUF_X1 U278 ( .A(n36), .Z(n302) );
  NOR2_X1 U279 ( .A1(n279), .A2(n324), .ZN(n303) );
  CLKBUF_X1 U280 ( .A(n70), .Z(n304) );
  NAND3_X1 U281 ( .A1(n309), .A2(n308), .A3(n307), .ZN(n305) );
  XOR2_X1 U282 ( .A(n85), .B(n84), .Z(n306) );
  XOR2_X1 U283 ( .A(n306), .B(n304), .Z(product[13]) );
  NAND2_X1 U284 ( .A1(n85), .A2(n84), .ZN(n307) );
  NAND2_X1 U285 ( .A1(n70), .A2(n85), .ZN(n308) );
  NAND2_X1 U286 ( .A1(n70), .A2(n84), .ZN(n309) );
  NAND3_X1 U287 ( .A1(n308), .A2(n307), .A3(n309), .ZN(n14) );
  NAND2_X1 U288 ( .A1(n141), .A2(n83), .ZN(n310) );
  NAND2_X1 U289 ( .A1(n305), .A2(n141), .ZN(n311) );
  NAND2_X1 U290 ( .A1(n83), .A2(n14), .ZN(n312) );
  XOR2_X1 U291 ( .A(n293), .B(a[4]), .Z(n314) );
  AOI21_X1 U292 ( .B1(n39), .B2(n47), .A(n40), .ZN(n315) );
  CLKBUF_X1 U293 ( .A(n29), .Z(n316) );
  XNOR2_X1 U294 ( .A(n236), .B(a[2]), .ZN(n317) );
  NAND2_X1 U295 ( .A1(n104), .A2(n109), .ZN(n318) );
  NAND2_X1 U296 ( .A1(n104), .A2(n106), .ZN(n319) );
  NAND2_X1 U297 ( .A1(n109), .A2(n106), .ZN(n320) );
  NAND3_X1 U298 ( .A1(n318), .A2(n319), .A3(n320), .ZN(n101) );
  BUF_X2 U299 ( .A(n216), .Z(n344) );
  CLKBUF_X1 U300 ( .A(n20), .Z(n321) );
  OAI22_X1 U301 ( .A1(n223), .A2(n192), .B1(n191), .B2(n342), .ZN(n322) );
  AOI21_X1 U302 ( .B1(n333), .B2(n55), .A(n52), .ZN(n323) );
  NOR2_X1 U303 ( .A1(n92), .A2(n95), .ZN(n324) );
  BUF_X2 U304 ( .A(n227), .Z(n342) );
  NOR2_X1 U305 ( .A1(n102), .A2(n107), .ZN(n325) );
  NAND2_X1 U306 ( .A1(n328), .A2(n294), .ZN(n326) );
  XNOR2_X1 U307 ( .A(n27), .B(n327), .ZN(product[11]) );
  AND2_X1 U308 ( .A1(n331), .A2(n26), .ZN(n327) );
  NOR2_X1 U309 ( .A1(n108), .A2(n113), .ZN(n44) );
  OR2_X1 U310 ( .A1(n88), .A2(n91), .ZN(n331) );
  NAND2_X1 U311 ( .A1(n281), .A2(n294), .ZN(n221) );
  XOR2_X1 U312 ( .A(n233), .B(a[6]), .Z(n328) );
  INV_X1 U313 ( .A(n279), .ZN(n74) );
  XOR2_X1 U314 ( .A(n37), .B(n329), .Z(product[9]) );
  AND2_X1 U315 ( .A1(n74), .A2(n302), .ZN(n329) );
  INV_X1 U316 ( .A(n302), .ZN(n34) );
  INV_X1 U317 ( .A(n26), .ZN(n24) );
  OAI21_X1 U318 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  NOR2_X1 U319 ( .A1(n102), .A2(n107), .ZN(n41) );
  AOI21_X1 U320 ( .B1(n330), .B2(n67), .A(n64), .ZN(n62) );
  INV_X1 U321 ( .A(n66), .ZN(n64) );
  NAND2_X1 U322 ( .A1(n332), .A2(n19), .ZN(n1) );
  XOR2_X1 U323 ( .A(n10), .B(n62), .Z(product[3]) );
  INV_X1 U324 ( .A(n60), .ZN(n80) );
  XOR2_X1 U325 ( .A(n9), .B(n58), .Z(product[4]) );
  NAND2_X1 U326 ( .A1(n79), .A2(n57), .ZN(n9) );
  INV_X1 U327 ( .A(n56), .ZN(n79) );
  XOR2_X1 U328 ( .A(n32), .B(n3), .Z(product[10]) );
  NAND2_X1 U329 ( .A1(n73), .A2(n31), .ZN(n3) );
  AOI21_X1 U330 ( .B1(n37), .B2(n74), .A(n34), .ZN(n32) );
  XOR2_X1 U331 ( .A(n46), .B(n6), .Z(product[7]) );
  NAND2_X1 U332 ( .A1(n76), .A2(n300), .ZN(n6) );
  INV_X1 U333 ( .A(n292), .ZN(n76) );
  NOR2_X1 U334 ( .A1(n101), .A2(n96), .ZN(n35) );
  XNOR2_X1 U335 ( .A(n43), .B(n5), .ZN(product[8]) );
  NAND2_X1 U336 ( .A1(n75), .A2(n42), .ZN(n5) );
  OAI21_X1 U337 ( .B1(n46), .B2(n292), .A(n300), .ZN(n43) );
  XNOR2_X1 U338 ( .A(n11), .B(n67), .ZN(product[2]) );
  NAND2_X1 U339 ( .A1(n330), .A2(n66), .ZN(n11) );
  XNOR2_X1 U340 ( .A(n8), .B(n55), .ZN(product[5]) );
  NAND2_X1 U341 ( .A1(n333), .A2(n54), .ZN(n8) );
  INV_X1 U342 ( .A(n59), .ZN(n58) );
  NAND2_X1 U343 ( .A1(n77), .A2(n49), .ZN(n7) );
  INV_X1 U344 ( .A(n48), .ZN(n77) );
  INV_X1 U345 ( .A(n19), .ZN(n17) );
  NOR2_X1 U346 ( .A1(n92), .A2(n95), .ZN(n30) );
  INV_X1 U347 ( .A(n69), .ZN(n67) );
  OR2_X1 U348 ( .A1(n171), .A2(n164), .ZN(n330) );
  NOR2_X1 U349 ( .A1(n122), .A2(n123), .ZN(n56) );
  NAND2_X1 U350 ( .A1(n108), .A2(n113), .ZN(n45) );
  NAND2_X1 U351 ( .A1(n114), .A2(n117), .ZN(n49) );
  NAND2_X1 U352 ( .A1(n88), .A2(n91), .ZN(n26) );
  NAND2_X1 U353 ( .A1(n87), .A2(n86), .ZN(n19) );
  NAND2_X1 U354 ( .A1(n124), .A2(n139), .ZN(n61) );
  NAND2_X1 U355 ( .A1(n122), .A2(n123), .ZN(n57) );
  NAND2_X1 U356 ( .A1(n92), .A2(n95), .ZN(n31) );
  OR2_X1 U357 ( .A1(n87), .A2(n86), .ZN(n332) );
  OR2_X1 U358 ( .A1(n344), .A2(n231), .ZN(n199) );
  AND2_X1 U359 ( .A1(n344), .A2(n129), .ZN(n156) );
  OAI22_X1 U360 ( .A1(n224), .A2(n204), .B1(n203), .B2(n244), .ZN(n169) );
  OAI22_X1 U361 ( .A1(n224), .A2(n203), .B1(n202), .B2(n244), .ZN(n168) );
  OAI22_X1 U362 ( .A1(n224), .A2(n202), .B1(n201), .B2(n244), .ZN(n167) );
  OR2_X1 U363 ( .A1(n344), .A2(n229), .ZN(n181) );
  AND2_X1 U364 ( .A1(n274), .A2(n69), .ZN(product[1]) );
  AND2_X1 U365 ( .A1(n344), .A2(n132), .ZN(n164) );
  OAI22_X1 U366 ( .A1(n224), .A2(n207), .B1(n206), .B2(n244), .ZN(n172) );
  OAI22_X1 U367 ( .A1(n224), .A2(n232), .B1(n208), .B2(n244), .ZN(n140) );
  OR2_X1 U368 ( .A1(n344), .A2(n232), .ZN(n208) );
  AND2_X1 U369 ( .A1(n344), .A2(n135), .ZN(product[0]) );
  INV_X1 U370 ( .A(n131), .ZN(n157) );
  NAND2_X1 U371 ( .A1(n171), .A2(n164), .ZN(n66) );
  OAI22_X1 U372 ( .A1(n224), .A2(n206), .B1(n205), .B2(n244), .ZN(n171) );
  INV_X1 U373 ( .A(n99), .ZN(n100) );
  NOR2_X1 U374 ( .A1(n124), .A2(n139), .ZN(n60) );
  OR2_X1 U375 ( .A1(n344), .A2(n230), .ZN(n190) );
  NAND2_X1 U376 ( .A1(n287), .A2(n226), .ZN(n222) );
  NAND2_X1 U377 ( .A1(n314), .A2(n301), .ZN(n337) );
  INV_X1 U378 ( .A(n125), .ZN(n141) );
  INV_X1 U379 ( .A(n83), .ZN(n84) );
  AND2_X1 U380 ( .A1(n344), .A2(n126), .ZN(n148) );
  OR2_X1 U381 ( .A1(n158), .A2(n146), .ZN(n105) );
  XNOR2_X1 U382 ( .A(n158), .B(n146), .ZN(n106) );
  INV_X1 U383 ( .A(n89), .ZN(n90) );
  INV_X1 U384 ( .A(n128), .ZN(n149) );
  INV_X1 U385 ( .A(n134), .ZN(n165) );
  AOI21_X1 U386 ( .B1(n37), .B2(n303), .A(n316), .ZN(n27) );
  NAND2_X1 U387 ( .A1(n80), .A2(n61), .ZN(n10) );
  OAI21_X1 U388 ( .B1(n60), .B2(n62), .A(n61), .ZN(n59) );
  XNOR2_X1 U389 ( .A(n235), .B(a[4]), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n235), .B(a[4]), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n235), .B(a[4]), .ZN(n226) );
  NAND2_X1 U392 ( .A1(n102), .A2(n107), .ZN(n42) );
  XNOR2_X1 U393 ( .A(n233), .B(b[6]), .ZN(n174) );
  XNOR2_X1 U394 ( .A(n233), .B(b[5]), .ZN(n175) );
  XNOR2_X1 U395 ( .A(n233), .B(b[4]), .ZN(n176) );
  XNOR2_X1 U396 ( .A(n233), .B(b[2]), .ZN(n178) );
  XNOR2_X1 U397 ( .A(n233), .B(b[3]), .ZN(n177) );
  XNOR2_X1 U398 ( .A(n344), .B(n233), .ZN(n180) );
  XNOR2_X1 U399 ( .A(n233), .B(b[1]), .ZN(n179) );
  INV_X1 U400 ( .A(n233), .ZN(n229) );
  NAND2_X1 U401 ( .A1(n96), .A2(n101), .ZN(n36) );
  NAND2_X2 U402 ( .A1(n220), .A2(n244), .ZN(n224) );
  NAND2_X1 U403 ( .A1(n219), .A2(n227), .ZN(n340) );
  NAND2_X1 U404 ( .A1(n313), .A2(n317), .ZN(n341) );
  NAND2_X1 U405 ( .A1(n313), .A2(n317), .ZN(n223) );
  XNOR2_X1 U406 ( .A(n236), .B(a[2]), .ZN(n227) );
  NAND2_X1 U407 ( .A1(n118), .A2(n121), .ZN(n54) );
  OAI22_X1 U408 ( .A1(n224), .A2(n205), .B1(n204), .B2(n244), .ZN(n170) );
  OAI21_X1 U409 ( .B1(n291), .B2(n323), .A(n49), .ZN(n343) );
  OAI21_X1 U410 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
  INV_X1 U411 ( .A(n324), .ZN(n73) );
  NOR2_X1 U412 ( .A1(n35), .A2(n324), .ZN(n28) );
  OAI21_X1 U413 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  XNOR2_X1 U414 ( .A(n236), .B(b[6]), .ZN(n201) );
  XNOR2_X1 U415 ( .A(n290), .B(b[5]), .ZN(n202) );
  XNOR2_X1 U416 ( .A(n290), .B(b[4]), .ZN(n203) );
  XNOR2_X1 U417 ( .A(n344), .B(n290), .ZN(n207) );
  INV_X1 U418 ( .A(n236), .ZN(n232) );
  INV_X1 U419 ( .A(n325), .ZN(n75) );
  NOR2_X1 U420 ( .A1(n325), .A2(n44), .ZN(n39) );
  OAI21_X1 U421 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  XNOR2_X1 U422 ( .A(n233), .B(b[7]), .ZN(n173) );
  OAI22_X1 U423 ( .A1(n224), .A2(n201), .B1(n200), .B2(n244), .ZN(n166) );
  OAI22_X1 U424 ( .A1(n200), .A2(n224), .B1(n200), .B2(n244), .ZN(n134) );
  AOI21_X1 U425 ( .B1(n333), .B2(n55), .A(n52), .ZN(n50) );
  NAND2_X1 U426 ( .A1(n28), .A2(n331), .ZN(n21) );
  AOI21_X1 U427 ( .B1(n29), .B2(n331), .A(n24), .ZN(n22) );
  OAI22_X1 U428 ( .A1(n173), .A2(n326), .B1(n173), .B2(n336), .ZN(n125) );
  OAI21_X1 U429 ( .B1(n38), .B2(n21), .A(n22), .ZN(n20) );
  OAI22_X1 U430 ( .A1(n326), .A2(n174), .B1(n173), .B2(n336), .ZN(n83) );
  OAI22_X1 U431 ( .A1(n326), .A2(n175), .B1(n174), .B2(n336), .ZN(n142) );
  OAI22_X1 U432 ( .A1(n326), .A2(n176), .B1(n175), .B2(n336), .ZN(n143) );
  OAI22_X1 U433 ( .A1(n326), .A2(n177), .B1(n176), .B2(n336), .ZN(n144) );
  INV_X1 U434 ( .A(n336), .ZN(n126) );
  OAI22_X1 U435 ( .A1(n326), .A2(n178), .B1(n177), .B2(n336), .ZN(n145) );
  OAI22_X1 U436 ( .A1(n326), .A2(n179), .B1(n178), .B2(n336), .ZN(n146) );
  OAI22_X1 U437 ( .A1(n221), .A2(n229), .B1(n181), .B2(n336), .ZN(n137) );
  OAI22_X1 U438 ( .A1(n180), .A2(n221), .B1(n179), .B2(n336), .ZN(n147) );
  XNOR2_X1 U439 ( .A(n236), .B(b[7]), .ZN(n200) );
  XNOR2_X1 U440 ( .A(n236), .B(b[1]), .ZN(n206) );
  XNOR2_X1 U441 ( .A(n290), .B(b[2]), .ZN(n205) );
  XNOR2_X1 U442 ( .A(n236), .B(b[3]), .ZN(n204) );
  INV_X1 U443 ( .A(n343), .ZN(n46) );
  AOI21_X1 U444 ( .B1(n47), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U445 ( .A1(n172), .A2(n140), .ZN(n69) );
  XOR2_X1 U446 ( .A(n7), .B(n323), .Z(product[6]) );
  OAI22_X1 U447 ( .A1(n182), .A2(n298), .B1(n182), .B2(n338), .ZN(n128) );
  OAI22_X1 U448 ( .A1(n337), .A2(n188), .B1(n187), .B2(n339), .ZN(n154) );
  OAI22_X1 U449 ( .A1(n298), .A2(n183), .B1(n182), .B2(n338), .ZN(n89) );
  OAI22_X1 U450 ( .A1(n337), .A2(n185), .B1(n184), .B2(n339), .ZN(n151) );
  OAI22_X1 U451 ( .A1(n289), .A2(n187), .B1(n186), .B2(n339), .ZN(n153) );
  OAI22_X1 U452 ( .A1(n289), .A2(n184), .B1(n183), .B2(n338), .ZN(n150) );
  OAI22_X1 U453 ( .A1(n337), .A2(n186), .B1(n185), .B2(n339), .ZN(n152) );
  INV_X1 U454 ( .A(n338), .ZN(n129) );
  XNOR2_X1 U455 ( .A(n280), .B(b[4]), .ZN(n194) );
  XNOR2_X1 U456 ( .A(n280), .B(b[5]), .ZN(n193) );
  XNOR2_X1 U457 ( .A(n280), .B(b[3]), .ZN(n195) );
  OAI22_X1 U458 ( .A1(n337), .A2(n230), .B1(n190), .B2(n339), .ZN(n138) );
  XNOR2_X1 U459 ( .A(n297), .B(b[2]), .ZN(n196) );
  INV_X1 U460 ( .A(n297), .ZN(n231) );
  XNOR2_X1 U461 ( .A(n235), .B(b[6]), .ZN(n192) );
  XNOR2_X1 U462 ( .A(n235), .B(b[7]), .ZN(n191) );
  XNOR2_X1 U463 ( .A(n344), .B(n297), .ZN(n198) );
  XNOR2_X1 U464 ( .A(n297), .B(b[1]), .ZN(n197) );
  XOR2_X1 U465 ( .A(n235), .B(a[2]), .Z(n219) );
  INV_X1 U466 ( .A(n15), .ZN(n70) );
  XNOR2_X1 U467 ( .A(n293), .B(b[7]), .ZN(n182) );
  XNOR2_X1 U468 ( .A(n293), .B(b[2]), .ZN(n187) );
  XNOR2_X1 U469 ( .A(n335), .B(b[5]), .ZN(n184) );
  XNOR2_X1 U470 ( .A(n293), .B(b[6]), .ZN(n183) );
  XNOR2_X1 U471 ( .A(n335), .B(b[3]), .ZN(n186) );
  XNOR2_X1 U472 ( .A(n293), .B(b[4]), .ZN(n185) );
  XNOR2_X1 U473 ( .A(n344), .B(n335), .ZN(n189) );
  INV_X1 U474 ( .A(n335), .ZN(n230) );
  XNOR2_X1 U475 ( .A(n293), .B(b[1]), .ZN(n188) );
  XOR2_X1 U476 ( .A(n335), .B(a[4]), .Z(n218) );
  XNOR2_X1 U477 ( .A(n321), .B(n1), .ZN(product[12]) );
  INV_X1 U478 ( .A(n315), .ZN(n37) );
  AOI21_X1 U479 ( .B1(n20), .B2(n332), .A(n17), .ZN(n15) );
  OAI22_X1 U480 ( .A1(n341), .A2(n193), .B1(n192), .B2(n296), .ZN(n158) );
  OAI22_X1 U481 ( .A1(n341), .A2(n195), .B1(n194), .B2(n296), .ZN(n160) );
  OAI22_X1 U482 ( .A1(n340), .A2(n194), .B1(n193), .B2(n342), .ZN(n159) );
  OAI22_X1 U483 ( .A1(n340), .A2(n196), .B1(n195), .B2(n342), .ZN(n161) );
  OAI22_X1 U484 ( .A1(n340), .A2(n231), .B1(n199), .B2(n342), .ZN(n139) );
  OAI22_X1 U485 ( .A1(n341), .A2(n197), .B1(n196), .B2(n296), .ZN(n162) );
  OAI22_X1 U486 ( .A1(n223), .A2(n192), .B1(n191), .B2(n342), .ZN(n99) );
  OAI22_X1 U487 ( .A1(n191), .A2(n340), .B1(n191), .B2(n342), .ZN(n131) );
  INV_X1 U488 ( .A(n342), .ZN(n132) );
  OAI22_X1 U489 ( .A1(n223), .A2(n198), .B1(n197), .B2(n296), .ZN(n163) );
  INV_X2 U490 ( .A(n135), .ZN(n244) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n54,
         n56, n57, n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  FA_X1 U6 ( .A(A[11]), .B(B[11]), .CI(n17), .CO(n16), .S(SUM[11]) );
  OR2_X1 U86 ( .A1(A[1]), .A2(B[1]), .ZN(n125) );
  OR2_X1 U87 ( .A1(A[0]), .A2(B[0]), .ZN(n126) );
  CLKBUF_X1 U88 ( .A(n25), .Z(n127) );
  CLKBUF_X1 U89 ( .A(n33), .Z(n128) );
  AOI21_X1 U90 ( .B1(n127), .B2(n139), .A(n22), .ZN(n129) );
  CLKBUF_X1 U91 ( .A(n41), .Z(n130) );
  AOI21_X1 U92 ( .B1(n133), .B2(n138), .A(n46), .ZN(n131) );
  AOI21_X1 U93 ( .B1(n125), .B2(n57), .A(n54), .ZN(n132) );
  CLKBUF_X1 U94 ( .A(n49), .Z(n133) );
  AOI21_X1 U95 ( .B1(n49), .B2(n138), .A(n46), .ZN(n44) );
  AOI21_X1 U96 ( .B1(n125), .B2(n57), .A(n54), .ZN(n52) );
  AOI21_X1 U97 ( .B1(n128), .B2(n140), .A(n30), .ZN(n134) );
  AOI21_X1 U98 ( .B1(n130), .B2(n137), .A(n38), .ZN(n135) );
  INV_X1 U99 ( .A(n24), .ZN(n22) );
  AOI21_X1 U100 ( .B1(n33), .B2(n140), .A(n30), .ZN(n28) );
  INV_X1 U101 ( .A(n32), .ZN(n30) );
  AOI21_X1 U102 ( .B1(n41), .B2(n137), .A(n38), .ZN(n36) );
  INV_X1 U103 ( .A(n40), .ZN(n38) );
  INV_X1 U104 ( .A(n56), .ZN(n54) );
  OAI21_X1 U105 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  INV_X1 U106 ( .A(n48), .ZN(n46) );
  NAND2_X1 U107 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U108 ( .A(n42), .ZN(n66) );
  NAND2_X1 U109 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U110 ( .A(n18), .ZN(n60) );
  NAND2_X1 U111 ( .A1(n138), .A2(n48), .ZN(n9) );
  NAND2_X1 U112 ( .A1(n139), .A2(n24), .ZN(n3) );
  XOR2_X1 U113 ( .A(n132), .B(n10), .Z(SUM[2]) );
  NAND2_X1 U114 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U115 ( .A(n50), .ZN(n68) );
  XOR2_X1 U116 ( .A(n135), .B(n6), .Z(SUM[6]) );
  NAND2_X1 U117 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U118 ( .A(n34), .ZN(n64) );
  XOR2_X1 U119 ( .A(n134), .B(n4), .Z(SUM[8]) );
  NAND2_X1 U120 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U121 ( .A(n26), .ZN(n62) );
  XNOR2_X1 U122 ( .A(n128), .B(n5), .ZN(SUM[7]) );
  NAND2_X1 U123 ( .A1(n140), .A2(n32), .ZN(n5) );
  XNOR2_X1 U124 ( .A(n130), .B(n7), .ZN(SUM[5]) );
  NAND2_X1 U125 ( .A1(n137), .A2(n40), .ZN(n7) );
  INV_X1 U126 ( .A(n59), .ZN(n57) );
  XNOR2_X1 U127 ( .A(n11), .B(n57), .ZN(SUM[1]) );
  NAND2_X1 U128 ( .A1(n125), .A2(n56), .ZN(n11) );
  XNOR2_X1 U129 ( .A(n13), .B(n136), .ZN(SUM[15]) );
  XNOR2_X1 U130 ( .A(B[15]), .B(A[15]), .ZN(n136) );
  NOR2_X1 U131 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  OR2_X1 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  OR2_X1 U133 ( .A1(A[3]), .A2(B[3]), .ZN(n138) );
  NOR2_X1 U134 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U135 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U136 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U137 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U138 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U140 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U141 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  NAND2_X1 U142 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  OR2_X1 U143 ( .A1(A[9]), .A2(B[9]), .ZN(n139) );
  OR2_X1 U144 ( .A1(A[7]), .A2(B[7]), .ZN(n140) );
  NAND2_X1 U145 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U146 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U147 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U148 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  AND2_X1 U149 ( .A1(n126), .A2(n59), .ZN(SUM[0]) );
  XNOR2_X1 U150 ( .A(n127), .B(n3), .ZN(SUM[9]) );
  AOI21_X1 U151 ( .B1(n25), .B2(n139), .A(n22), .ZN(n20) );
  OAI21_X1 U152 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U153 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  XOR2_X1 U154 ( .A(n131), .B(n8), .Z(SUM[4]) );
  XNOR2_X1 U155 ( .A(n133), .B(n9), .ZN(SUM[3]) );
  XOR2_X1 U156 ( .A(n129), .B(n2), .Z(SUM[10]) );
  NAND2_X1 U157 ( .A1(A[0]), .A2(B[0]), .ZN(n59) );
  NAND2_X1 U158 ( .A1(A[1]), .A2(B[1]), .ZN(n56) );
  OAI21_X1 U159 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X1 U160 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
endmodule


module add_layer_WIDTH16_6 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_6_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n54,
         n56, n57, n59, n60, n62, n64, n66, n68, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n14), .CO(n13), .S(SUM[14]) );
  FA_X1 U4 ( .A(A[13]), .B(B[13]), .CI(n15), .CO(n14), .S(SUM[13]) );
  FA_X1 U5 ( .A(A[12]), .B(B[12]), .CI(n16), .CO(n15), .S(SUM[12]) );
  AOI21_X1 U86 ( .B1(n49), .B2(n141), .A(n46), .ZN(n44) );
  OR2_X1 U87 ( .A1(A[0]), .A2(B[0]), .ZN(n125) );
  AOI21_X1 U88 ( .B1(n138), .B2(n57), .A(n54), .ZN(n126) );
  AOI21_X1 U89 ( .B1(n138), .B2(n57), .A(n54), .ZN(n52) );
  XOR2_X1 U90 ( .A(A[11]), .B(B[11]), .Z(n127) );
  XOR2_X1 U91 ( .A(n17), .B(n127), .Z(SUM[11]) );
  NAND2_X1 U92 ( .A1(n17), .A2(A[11]), .ZN(n128) );
  NAND2_X1 U93 ( .A1(n17), .A2(B[11]), .ZN(n129) );
  NAND2_X1 U94 ( .A1(A[11]), .A2(B[11]), .ZN(n130) );
  NAND3_X1 U95 ( .A1(n128), .A2(n129), .A3(n130), .ZN(n16) );
  CLKBUF_X1 U96 ( .A(n33), .Z(n131) );
  CLKBUF_X1 U97 ( .A(n49), .Z(n132) );
  CLKBUF_X1 U98 ( .A(n41), .Z(n133) );
  CLKBUF_X1 U99 ( .A(n25), .Z(n134) );
  AOI21_X1 U100 ( .B1(n133), .B2(n140), .A(n38), .ZN(n135) );
  AOI21_X1 U101 ( .B1(n134), .B2(n142), .A(n22), .ZN(n136) );
  AOI21_X1 U102 ( .B1(n131), .B2(n143), .A(n30), .ZN(n137) );
  INV_X1 U103 ( .A(n24), .ZN(n22) );
  AOI21_X1 U104 ( .B1(n33), .B2(n143), .A(n30), .ZN(n28) );
  INV_X1 U105 ( .A(n32), .ZN(n30) );
  INV_X1 U106 ( .A(n48), .ZN(n46) );
  AOI21_X1 U107 ( .B1(n41), .B2(n140), .A(n38), .ZN(n36) );
  INV_X1 U108 ( .A(n40), .ZN(n38) );
  NAND2_X1 U109 ( .A1(n60), .A2(n19), .ZN(n2) );
  INV_X1 U110 ( .A(n18), .ZN(n60) );
  NAND2_X1 U111 ( .A1(n66), .A2(n43), .ZN(n8) );
  INV_X1 U112 ( .A(n42), .ZN(n66) );
  NAND2_X1 U113 ( .A1(n64), .A2(n35), .ZN(n6) );
  INV_X1 U114 ( .A(n34), .ZN(n64) );
  NAND2_X1 U115 ( .A1(n62), .A2(n27), .ZN(n4) );
  INV_X1 U116 ( .A(n26), .ZN(n62) );
  INV_X1 U117 ( .A(n56), .ZN(n54) );
  NAND2_X1 U118 ( .A1(n143), .A2(n32), .ZN(n5) );
  NAND2_X1 U119 ( .A1(n142), .A2(n24), .ZN(n3) );
  INV_X1 U120 ( .A(n59), .ZN(n57) );
  XNOR2_X1 U121 ( .A(n132), .B(n9), .ZN(SUM[3]) );
  NAND2_X1 U122 ( .A1(n141), .A2(n48), .ZN(n9) );
  XNOR2_X1 U123 ( .A(n133), .B(n7), .ZN(SUM[5]) );
  NAND2_X1 U124 ( .A1(n140), .A2(n40), .ZN(n7) );
  XNOR2_X1 U125 ( .A(n11), .B(n57), .ZN(SUM[1]) );
  NAND2_X1 U126 ( .A1(n138), .A2(n56), .ZN(n11) );
  NAND2_X1 U127 ( .A1(n68), .A2(n51), .ZN(n10) );
  INV_X1 U128 ( .A(n50), .ZN(n68) );
  OR2_X1 U129 ( .A1(A[1]), .A2(B[1]), .ZN(n138) );
  XNOR2_X1 U130 ( .A(n13), .B(n139), .ZN(SUM[15]) );
  XNOR2_X1 U131 ( .A(B[15]), .B(A[15]), .ZN(n139) );
  OR2_X1 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n140) );
  OR2_X1 U133 ( .A1(A[3]), .A2(B[3]), .ZN(n141) );
  NOR2_X1 U134 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  NOR2_X1 U135 ( .A1(A[6]), .A2(B[6]), .ZN(n34) );
  NOR2_X1 U136 ( .A1(A[2]), .A2(B[2]), .ZN(n50) );
  NOR2_X1 U137 ( .A1(A[8]), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U138 ( .A1(A[10]), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(n32) );
  NAND2_X1 U140 ( .A1(A[5]), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U141 ( .A1(A[3]), .A2(B[3]), .ZN(n48) );
  NAND2_X1 U142 ( .A1(A[9]), .A2(B[9]), .ZN(n24) );
  OR2_X1 U143 ( .A1(A[9]), .A2(B[9]), .ZN(n142) );
  OR2_X1 U144 ( .A1(A[7]), .A2(B[7]), .ZN(n143) );
  NAND2_X1 U145 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  NAND2_X1 U146 ( .A1(A[6]), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U147 ( .A1(A[2]), .A2(B[2]), .ZN(n51) );
  NAND2_X1 U148 ( .A1(A[8]), .A2(B[8]), .ZN(n27) );
  NAND2_X1 U149 ( .A1(A[10]), .A2(B[10]), .ZN(n19) );
  AND2_X1 U150 ( .A1(n125), .A2(n59), .ZN(SUM[0]) );
  XOR2_X1 U151 ( .A(n135), .B(n6), .Z(SUM[6]) );
  XOR2_X1 U152 ( .A(n44), .B(n8), .Z(SUM[4]) );
  OAI21_X1 U153 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  NAND2_X1 U154 ( .A1(A[0]), .A2(B[0]), .ZN(n59) );
  XNOR2_X1 U155 ( .A(n131), .B(n5), .ZN(SUM[7]) );
  OAI21_X1 U156 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U157 ( .A(n134), .B(n3), .ZN(SUM[9]) );
  XOR2_X1 U158 ( .A(n126), .B(n10), .Z(SUM[2]) );
  XOR2_X1 U159 ( .A(n136), .B(n2), .Z(SUM[10]) );
  AOI21_X1 U160 ( .B1(n25), .B2(n142), .A(n22), .ZN(n20) );
  OAI21_X1 U161 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  NAND2_X1 U162 ( .A1(A[1]), .A2(B[1]), .ZN(n56) );
  OAI21_X1 U163 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U164 ( .B1(n20), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U165 ( .A(n137), .B(n4), .Z(SUM[8]) );
endmodule


module add_layer_WIDTH16_5 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_5_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n19, n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37,
         n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55,
         n56, n57, n61, n64, n65, n67, n69, n71, n73, n75, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n162, n163, n164;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n15), .CO(n14), .S(SUM[14]) );
  INV_X1 U94 ( .A(n144), .ZN(n64) );
  OR2_X1 U95 ( .A1(A[0]), .A2(B[0]), .ZN(n132) );
  CLKBUF_X1 U96 ( .A(n157), .Z(n133) );
  OR2_X1 U97 ( .A1(B[1]), .A2(A[1]), .ZN(n157) );
  CLKBUF_X1 U98 ( .A(n54), .Z(n134) );
  AND2_X1 U99 ( .A1(A[1]), .A2(B[1]), .ZN(n154) );
  INV_X1 U100 ( .A(n154), .ZN(n61) );
  CLKBUF_X1 U101 ( .A(n138), .Z(n135) );
  AOI21_X1 U102 ( .B1(n134), .B2(n159), .A(n51), .ZN(n136) );
  AOI21_X1 U103 ( .B1(n54), .B2(n159), .A(n51), .ZN(n49) );
  CLKBUF_X1 U104 ( .A(n30), .Z(n137) );
  NAND3_X1 U105 ( .A1(n148), .A2(n147), .A3(n146), .ZN(n138) );
  AOI21_X1 U106 ( .B1(n137), .B2(n162), .A(n27), .ZN(n139) );
  CLKBUF_X1 U107 ( .A(n46), .Z(n140) );
  CLKBUF_X1 U108 ( .A(n22), .Z(n141) );
  AOI21_X1 U109 ( .B1(n30), .B2(n162), .A(n27), .ZN(n25) );
  CLKBUF_X1 U110 ( .A(n65), .Z(n142) );
  AOI21_X1 U111 ( .B1(n140), .B2(n160), .A(n43), .ZN(n143) );
  AOI21_X1 U112 ( .B1(n46), .B2(n160), .A(n43), .ZN(n41) );
  AND2_X2 U113 ( .A1(A[0]), .A2(B[0]), .ZN(n144) );
  XOR2_X1 U114 ( .A(A[12]), .B(B[12]), .Z(n145) );
  XOR2_X1 U115 ( .A(n145), .B(n142), .Z(SUM[12]) );
  NAND2_X1 U116 ( .A1(A[12]), .A2(B[12]), .ZN(n146) );
  NAND2_X1 U117 ( .A1(n65), .A2(A[12]), .ZN(n147) );
  NAND2_X1 U118 ( .A1(n65), .A2(B[12]), .ZN(n148) );
  NAND3_X1 U119 ( .A1(n147), .A2(n146), .A3(n148), .ZN(n16) );
  XOR2_X1 U120 ( .A(A[13]), .B(B[13]), .Z(n149) );
  XOR2_X1 U121 ( .A(n149), .B(n135), .Z(SUM[13]) );
  NAND2_X1 U122 ( .A1(A[13]), .A2(B[13]), .ZN(n150) );
  NAND2_X1 U123 ( .A1(n138), .A2(A[13]), .ZN(n151) );
  NAND2_X1 U124 ( .A1(B[13]), .A2(n16), .ZN(n152) );
  NAND3_X1 U125 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n15) );
  CLKBUF_X1 U126 ( .A(n38), .Z(n153) );
  AOI21_X1 U127 ( .B1(n38), .B2(n163), .A(n35), .ZN(n155) );
  AOI21_X1 U128 ( .B1(n157), .B2(n144), .A(n154), .ZN(n156) );
  INV_X1 U129 ( .A(n29), .ZN(n27) );
  INV_X1 U130 ( .A(n37), .ZN(n35) );
  INV_X1 U131 ( .A(n53), .ZN(n51) );
  INV_X1 U132 ( .A(n45), .ZN(n43) );
  AOI21_X1 U133 ( .B1(n133), .B2(n144), .A(n154), .ZN(n57) );
  NAND2_X1 U134 ( .A1(n67), .A2(n24), .ZN(n3) );
  INV_X1 U135 ( .A(n23), .ZN(n67) );
  NAND2_X1 U136 ( .A1(n73), .A2(n48), .ZN(n9) );
  INV_X1 U137 ( .A(n47), .ZN(n73) );
  NAND2_X1 U138 ( .A1(n71), .A2(n40), .ZN(n7) );
  INV_X1 U139 ( .A(n39), .ZN(n71) );
  NAND2_X1 U140 ( .A1(n69), .A2(n32), .ZN(n5) );
  INV_X1 U141 ( .A(n31), .ZN(n69) );
  NAND2_X1 U142 ( .A1(n164), .A2(n21), .ZN(n2) );
  NAND2_X1 U143 ( .A1(n162), .A2(n29), .ZN(n4) );
  NAND2_X1 U144 ( .A1(n159), .A2(n53), .ZN(n10) );
  NAND2_X1 U145 ( .A1(n160), .A2(n45), .ZN(n8) );
  NAND2_X1 U146 ( .A1(n163), .A2(n37), .ZN(n6) );
  NAND2_X1 U147 ( .A1(n75), .A2(n56), .ZN(n11) );
  INV_X1 U148 ( .A(n55), .ZN(n75) );
  XNOR2_X1 U149 ( .A(n14), .B(n158), .ZN(SUM[15]) );
  XNOR2_X1 U150 ( .A(B[15]), .B(A[15]), .ZN(n158) );
  INV_X1 U151 ( .A(n21), .ZN(n19) );
  OR2_X1 U152 ( .A1(A[3]), .A2(B[3]), .ZN(n159) );
  OR2_X1 U153 ( .A1(A[5]), .A2(B[5]), .ZN(n160) );
  NOR2_X1 U154 ( .A1(A[8]), .A2(B[8]), .ZN(n31) );
  NOR2_X1 U155 ( .A1(A[6]), .A2(B[6]), .ZN(n39) );
  NOR2_X1 U156 ( .A1(A[2]), .A2(B[2]), .ZN(n55) );
  NOR2_X1 U157 ( .A1(A[4]), .A2(B[4]), .ZN(n47) );
  NOR2_X1 U158 ( .A1(A[10]), .A2(B[10]), .ZN(n23) );
  AND2_X1 U159 ( .A1(n132), .A2(n64), .ZN(SUM[0]) );
  NAND2_X1 U160 ( .A1(A[9]), .A2(B[9]), .ZN(n29) );
  NAND2_X1 U161 ( .A1(A[7]), .A2(B[7]), .ZN(n37) );
  NAND2_X1 U162 ( .A1(A[3]), .A2(B[3]), .ZN(n53) );
  NAND2_X1 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n45) );
  NAND2_X1 U164 ( .A1(A[11]), .A2(B[11]), .ZN(n21) );
  OR2_X1 U165 ( .A1(A[9]), .A2(B[9]), .ZN(n162) );
  OR2_X1 U166 ( .A1(A[7]), .A2(B[7]), .ZN(n163) );
  OR2_X1 U167 ( .A1(A[11]), .A2(B[11]), .ZN(n164) );
  NAND2_X1 U168 ( .A1(A[8]), .A2(B[8]), .ZN(n32) );
  NAND2_X1 U169 ( .A1(A[6]), .A2(B[6]), .ZN(n40) );
  NAND2_X1 U170 ( .A1(A[2]), .A2(B[2]), .ZN(n56) );
  NAND2_X1 U171 ( .A1(A[4]), .A2(B[4]), .ZN(n48) );
  NAND2_X1 U172 ( .A1(A[10]), .A2(B[10]), .ZN(n24) );
  XNOR2_X1 U173 ( .A(n12), .B(n144), .ZN(SUM[1]) );
  NAND2_X1 U174 ( .A1(n133), .A2(n61), .ZN(n12) );
  XNOR2_X1 U175 ( .A(n141), .B(n2), .ZN(SUM[11]) );
  XNOR2_X1 U176 ( .A(n137), .B(n4), .ZN(SUM[9]) );
  XNOR2_X1 U177 ( .A(n153), .B(n6), .ZN(SUM[7]) );
  XOR2_X1 U178 ( .A(n33), .B(n5), .Z(SUM[8]) );
  INV_X1 U179 ( .A(n17), .ZN(n65) );
  AOI21_X1 U180 ( .B1(n153), .B2(n163), .A(n35), .ZN(n33) );
  OAI21_X1 U181 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U182 ( .B1(n155), .B2(n31), .A(n32), .ZN(n30) );
  AOI21_X1 U183 ( .B1(n22), .B2(n164), .A(n19), .ZN(n17) );
  XOR2_X1 U184 ( .A(n143), .B(n7), .Z(SUM[6]) );
  XOR2_X1 U185 ( .A(n139), .B(n3), .Z(SUM[10]) );
  OAI21_X1 U186 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
  XNOR2_X1 U187 ( .A(n140), .B(n8), .ZN(SUM[5]) );
  OAI21_X1 U188 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  XOR2_X1 U189 ( .A(n136), .B(n9), .Z(SUM[4]) );
  XNOR2_X1 U190 ( .A(n134), .B(n10), .ZN(SUM[3]) );
  OAI21_X1 U191 ( .B1(n156), .B2(n55), .A(n56), .ZN(n54) );
  XOR2_X1 U192 ( .A(n57), .B(n11), .Z(SUM[2]) );
endmodule


module add_layer_WIDTH16_1 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_1_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_1 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_1 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_1 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_6 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_5 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_1 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_1 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4 \genblk1[0].mult  ( .clk(clk), .ia(
        {\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3 \genblk1[1].mult  ( .clk(clk), .ia(
        {\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2 \genblk1[2].mult  ( .clk(clk), .ia(
        {\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1 \genblk1[3].mult  ( .clk(clk), .ia(
        {\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_1 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module data_path_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_DELAY2 ( clk, 
        en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay, of_a, 
        of_x, of_y, of_delay, data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay;
  output of_a, of_x, of_y, of_delay;
  wire   N24, N25, \a[15][7] , \a[15][6] , \a[15][5] , \a[15][4] , \a[15][3] ,
         \a[15][2] , \a[15][1] , \a[15][0] , \a[14][7] , \a[14][6] ,
         \a[14][5] , \a[14][4] , \a[14][3] , \a[14][2] , \a[14][0] ,
         \a[13][7] , \a[13][6] , \a[13][5] , \a[13][4] , \a[13][3] ,
         \a[13][2] , \a[13][1] , \a[13][0] , \a[12][7] , \a[12][6] ,
         \a[12][5] , \a[12][4] , \a[12][2] , \a[12][1] , \a[12][0] ,
         \a[11][7] , \a[11][6] , \a[11][5] , \a[11][4] , \a[11][3] ,
         \a[11][2] , \a[11][1] , \a[11][0] , \a[10][7] , \a[10][6] ,
         \a[10][5] , \a[10][4] , \a[10][3] , \a[10][2] , \a[10][1] ,
         \a[10][0] , \a[9][7] , \a[9][6] , \a[9][5] , \a[9][4] , \a[9][3] ,
         \a[9][2] , \a[9][1] , \a[9][0] , \a[8][7] , \a[8][6] , \a[8][5] ,
         \a[8][4] , \a[8][3] , \a[8][2] , \a[8][1] , \a[8][0] , \a[7][7] ,
         \a[7][6] , \a[7][5] , \a[7][4] , \a[7][3] , \a[7][2] , \a[7][1] ,
         \a[7][0] , \a[6][7] , \a[6][6] , \a[6][5] , \a[6][4] , \a[6][3] ,
         \a[6][2] , \a[6][0] , \a[5][7] , \a[5][6] , \a[5][5] , \a[5][4] ,
         \a[5][3] , \a[5][2] , \a[5][0] , \a[4][7] , \a[4][6] , \a[4][5] ,
         \a[4][4] , \a[4][2] , \a[4][1] , \a[4][0] , \a[3][7] , \a[3][6] ,
         \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , \a[3][0] ,
         \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] ,
         \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] ,
         \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , \a[0][6] ,
         \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , \a[0][0] ,
         \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , \x[3][2] ,
         \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] ,
         \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , \x[1][7] , \x[1][6] ,
         \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] ,
         \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , \x[0][2] ,
         \x[0][1] , \x[0][0] , \y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] ,
         \y[3][11] , \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] ,
         \y[3][5] , \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] ,
         \y[2][15] , \y[2][14] , \y[2][13] , \y[2][12] , \y[2][11] ,
         \y[2][10] , \y[2][9] , \y[2][8] , \y[2][7] , \y[2][6] , \y[2][5] ,
         \y[2][4] , \y[2][3] , \y[2][2] , \y[2][1] , \y[2][0] , \y[1][15] ,
         \y[1][14] , \y[1][13] , \y[1][12] , \y[1][11] , \y[1][10] , \y[1][9] ,
         \y[1][8] , \y[1][7] , \y[1][6] , \y[1][5] , \y[1][4] , \y[1][3] ,
         \y[1][2] , \y[1][1] , \y[1][0] , \y[0][15] , \y[0][14] , \y[0][13] ,
         \y[0][12] , \y[0][11] , \y[0][10] , \y[0][9] , \y[0][8] , \y[0][7] ,
         \y[0][6] , \y[0][5] , \y[0][4] , \y[0][3] , \y[0][2] , \y[0][1] ,
         \y[0][0] , N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N89, N91, N92, N96, N97, N101, N102, N108, N109,
         N110, N114, N115, N116, n9, n10, n12, n15, n16, n19, n20, n21, n32,
         n38, n39, n40, n41, n47, n48, n49, n50, n51, n52, n58, n59, n60, n61,
         n62, n68, n69, n70, n71, n72, n78, n79, n80, n81, n82, n88, n89, n90,
         n91, n97, n98, n99, n100, n101, n102, n103, n107, n108, n109, n110,
         n111, n112, n116, n117, n118, n119, n120, n121, n125, n126, n127,
         n128, n129, n130, n134, n135, n136, n137, n143, n144, n145, n146,
         n152, n153, n154, n155, n156, n162, n163, n164, n165, n171, n172,
         n173, n174, n175, n181, n182, n183, n184, n185, n191, n192, n193,
         n194, n200, n201, n202, n203, n209, n210, n211, n212, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n1, n2, n3, n4, n5, n6, n7, n8, n11, n13, n14, n17, n18, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37,
         n42, n43, n44, n45, n46, n53, n54, n55, n56, n57, n63, n64, n65, n66,
         n67, n73, n74, n75, n76, n77, n83, n84, n85, n86, n87, n92, n93, n94,
         n95, n96, n104, n105, n106, n113, n114, n115, n122, n123, n124, n131,
         n132, n133, n138, n139, n140, n141, n142, n147, n148, n149, n150,
         n151, n157, n158, n159, n160, n161, n166, n167, n168, n169, n170,
         n176, n177, n178, n179, n180, n186, n187, n188, n189, n190, n195,
         n196, n197, n198, n199, n204, n205, n206, n207, n208, n213, n214,
         n215, n216, n217, n230, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443;
  wire   [3:0] addr_a;
  wire   [1:0] addr_x;
  wire   [3:0] delay_timer;
  assign of_a = N114;
  assign of_x = N115;
  assign of_y = N116;

  DFF_X1 \data_out_reg[15]  ( .D(N68), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N69), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N70), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N71), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N72), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N73), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N74), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N75), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N76), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N77), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N78), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N79), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N80), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N81), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N82), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N83), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \addr_a_reg[0]  ( .D(N89), .CK(clk), .Q(addr_a[0]) );
  DFF_X1 \addr_a_reg[1]  ( .D(n435), .CK(clk), .Q(addr_a[1]), .QN(n12) );
  DFF_X1 \addr_a_reg[2]  ( .D(N91), .CK(clk), .Q(addr_a[2]), .QN(n10) );
  DFF_X1 \addr_a_reg[3]  ( .D(N92), .CK(clk), .Q(addr_a[3]), .QN(n9) );
  DFF_X1 \a_reg[3][6]  ( .D(n356), .CK(clk), .Q(\a[3][6] ) );
  DFF_X1 \a_reg[3][4]  ( .D(n358), .CK(clk), .Q(\a[3][4] ) );
  DFF_X1 \a_reg[3][2]  ( .D(n360), .CK(clk), .Q(\a[3][2] ) );
  DFF_X1 \a_reg[3][0]  ( .D(n362), .CK(clk), .Q(\a[3][0] ) );
  DFF_X1 \a_reg[2][6]  ( .D(n364), .CK(clk), .Q(\a[2][6] ) );
  DFF_X1 \a_reg[2][4]  ( .D(n366), .CK(clk), .Q(\a[2][4] ) );
  DFF_X1 \a_reg[2][0]  ( .D(n370), .CK(clk), .Q(\a[2][0] ) );
  DFF_X1 \a_reg[1][6]  ( .D(n372), .CK(clk), .Q(\a[1][6] ) );
  DFF_X1 \a_reg[1][4]  ( .D(n374), .CK(clk), .Q(\a[1][4] ) );
  DFF_X1 \a_reg[1][2]  ( .D(n376), .CK(clk), .Q(\a[1][2] ) );
  DFF_X1 \a_reg[1][0]  ( .D(n378), .CK(clk), .Q(\a[1][0] ) );
  DFF_X1 \a_reg[0][6]  ( .D(n380), .CK(clk), .Q(\a[0][6] ) );
  DFF_X1 \a_reg[0][4]  ( .D(n382), .CK(clk), .Q(\a[0][4] ) );
  DFF_X1 \a_reg[0][2]  ( .D(n384), .CK(clk), .Q(\a[0][2] ) );
  DFF_X1 \a_reg[0][0]  ( .D(n386), .CK(clk), .Q(\a[0][0] ) );
  DFF_X1 \a_reg[11][6]  ( .D(n292), .CK(clk), .Q(\a[11][6] ) );
  DFF_X1 \a_reg[11][4]  ( .D(n294), .CK(clk), .Q(\a[11][4] ) );
  DFF_X1 \a_reg[11][2]  ( .D(n296), .CK(clk), .Q(\a[11][2] ) );
  DFF_X1 \a_reg[10][7]  ( .D(n299), .CK(clk), .Q(\a[10][7] ), .QN(n45) );
  DFF_X1 \a_reg[10][6]  ( .D(n300), .CK(clk), .Q(\a[10][6] ) );
  DFF_X1 \a_reg[10][4]  ( .D(n302), .CK(clk), .Q(\a[10][4] ) );
  DFF_X1 \a_reg[10][2]  ( .D(n304), .CK(clk), .Q(\a[10][2] ) );
  DFF_X1 \a_reg[10][0]  ( .D(n306), .CK(clk), .Q(\a[10][0] ) );
  DFF_X1 \a_reg[9][6]  ( .D(n308), .CK(clk), .Q(\a[9][6] ) );
  DFF_X1 \a_reg[9][4]  ( .D(n310), .CK(clk), .Q(\a[9][4] ) );
  DFF_X1 \a_reg[8][6]  ( .D(n316), .CK(clk), .Q(\a[8][6] ) );
  DFF_X1 \a_reg[8][4]  ( .D(n318), .CK(clk), .Q(\a[8][4] ) );
  DFF_X1 \a_reg[8][2]  ( .D(n320), .CK(clk), .Q(\a[8][2] ) );
  DFF_X1 \a_reg[8][0]  ( .D(n322), .CK(clk), .Q(\a[8][0] ) );
  DFF_X1 \a_reg[14][6]  ( .D(n268), .CK(clk), .Q(\a[14][6] ) );
  DFF_X1 \a_reg[14][4]  ( .D(n270), .CK(clk), .Q(\a[14][4] ) );
  DFF_X1 \a_reg[14][0]  ( .D(n274), .CK(clk), .Q(\a[14][0] ) );
  DFF_X1 \a_reg[13][6]  ( .D(n276), .CK(clk), .Q(\a[13][6] ) );
  DFF_X1 \a_reg[13][4]  ( .D(n278), .CK(clk), .Q(\a[13][4] ) );
  DFF_X1 \a_reg[13][2]  ( .D(n280), .CK(clk), .Q(\a[13][2] ) );
  DFF_X1 \a_reg[13][0]  ( .D(n282), .CK(clk), .Q(\a[13][0] ) );
  DFF_X1 \a_reg[12][7]  ( .D(n283), .CK(clk), .Q(\a[12][7] ) );
  DFF_X1 \a_reg[12][6]  ( .D(n284), .CK(clk), .Q(\a[12][6] ) );
  DFF_X1 \a_reg[12][4]  ( .D(n286), .CK(clk), .Q(\a[12][4] ) );
  DFF_X1 \a_reg[12][2]  ( .D(n288), .CK(clk), .Q(\a[12][2] ) );
  DFF_X1 \a_reg[12][0]  ( .D(n290), .CK(clk), .Q(\a[12][0] ) );
  DFF_X1 \a_reg[5][7]  ( .D(n339), .CK(clk), .Q(\a[5][7] ), .QN(n73) );
  DFF_X1 \a_reg[5][6]  ( .D(n340), .CK(clk), .Q(\a[5][6] ) );
  DFF_X1 \a_reg[5][4]  ( .D(n342), .CK(clk), .Q(\a[5][4] ) );
  DFF_X1 \a_reg[5][2]  ( .D(n344), .CK(clk), .Q(\a[5][2] ) );
  DFF_X1 \a_reg[5][0]  ( .D(n346), .CK(clk), .Q(\a[5][0] ) );
  DFF_X1 \a_reg[4][6]  ( .D(n348), .CK(clk), .Q(\a[4][6] ) );
  DFF_X1 \a_reg[4][2]  ( .D(n352), .CK(clk), .Q(\a[4][2] ) );
  DFF_X1 \a_reg[4][0]  ( .D(n354), .CK(clk), .Q(\a[4][0] ) );
  DFF_X1 \a_reg[7][7]  ( .D(n323), .CK(clk), .Q(\a[7][7] ) );
  DFF_X1 \a_reg[7][2]  ( .D(n328), .CK(clk), .Q(\a[7][2] ) );
  DFF_X1 \a_reg[7][0]  ( .D(n330), .CK(clk), .Q(\a[7][0] ) );
  DFF_X1 \a_reg[6][4]  ( .D(n334), .CK(clk), .Q(\a[6][4] ) );
  DFF_X1 \a_reg[6][2]  ( .D(n336), .CK(clk), .Q(\a[6][2] ) );
  DFF_X1 \a_reg[6][0]  ( .D(n338), .CK(clk), .Q(\a[6][0] ) );
  DFF_X1 \a_reg[6][6]  ( .D(n332), .CK(clk), .Q(\a[6][6] ) );
  DFF_X1 \a_reg[15][6]  ( .D(n260), .CK(clk), .Q(\a[15][6] ) );
  DFF_X1 \a_reg[15][4]  ( .D(n262), .CK(clk), .Q(\a[15][4] ) );
  DFF_X1 \a_reg[15][2]  ( .D(n264), .CK(clk), .Q(\a[15][2] ) );
  DFF_X1 \a_reg[15][0]  ( .D(n266), .CK(clk), .Q(\a[15][0] ) );
  DFF_X1 \addr_x_reg[0]  ( .D(N96), .CK(clk), .Q(addr_x[0]), .QN(n16) );
  DFF_X1 \addr_x_reg[1]  ( .D(N97), .CK(clk), .Q(addr_x[1]), .QN(n15) );
  DFF_X1 \x_reg[2][5]  ( .D(n237), .CK(clk), .Q(\x[2][5] ) );
  DFF_X1 \x_reg[2][0]  ( .D(n242), .CK(clk), .Q(\x[2][0] ) );
  DFF_X1 \x_reg[0][7]  ( .D(n251), .CK(clk), .Q(\x[0][7] ), .QN(n43) );
  DFF_X1 \x_reg[0][3]  ( .D(n255), .CK(clk), .Q(\x[0][3] ), .QN(n35) );
  DFF_X1 \x_reg[0][0]  ( .D(n258), .CK(clk), .Q(\x[0][0] ) );
  DFF_X1 \x_reg[1][0]  ( .D(n250), .CK(clk), .Q(\x[1][0] ) );
  DFF_X1 \x_reg[3][7]  ( .D(n426), .CK(clk), .Q(\x[3][7] ), .QN(n30) );
  DFF_X1 \x_reg[3][5]  ( .D(n428), .CK(clk), .Q(\x[3][5] ) );
  DFF_X1 \x_reg[3][0]  ( .D(n433), .CK(clk), .Q(\x[3][0] ) );
  DFF_X1 \addr_y_reg[1]  ( .D(N102), .CK(clk), .Q(N25), .QN(n3) );
  DFF_X1 \delay_timer_reg[0]  ( .D(N108), .CK(clk), .Q(delay_timer[0]), .QN(
        n21) );
  DFF_X1 \delay_timer_reg[1]  ( .D(N109), .CK(clk), .Q(delay_timer[1]), .QN(
        n20) );
  DFF_X1 \delay_timer_reg[2]  ( .D(N110), .CK(clk), .Q(delay_timer[2]), .QN(
        n19) );
  DFF_X1 \delay_timer_reg[3]  ( .D(n437), .CK(clk), .Q(delay_timer[3]) );
  NAND3_X1 U394 ( .A1(delay_timer[0]), .A2(n438), .A3(delay_timer[1]), .ZN(
        n231) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_0 \genblk1[0].element  ( 
        .clk(clk), .a({n115, \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , 
        \a[3][2] , \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , n133, \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , n131, \a[1][6] , \a[1][5] , 
        \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .x({\x[3][7] , \x[3][6] , n214, \x[3][4] , \x[3][3] , 
        \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , n29, n215, \x[2][4] , 
        \x[2][3] , \x[2][2] , n87, \x[2][0] , \x[1][7] , \x[1][6] , \x[1][5] , 
        n6, \x[1][3] , \x[1][2] , n85, \x[1][0] , n44, \x[0][6] , n217, 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .y({
        \y[0][15] , \y[0][14] , \y[0][13] , \y[0][12] , \y[0][11] , \y[0][10] , 
        \y[0][9] , \y[0][8] , \y[0][7] , \y[0][6] , \y[0][5] , \y[0][4] , 
        \y[0][3] , \y[0][2] , \y[0][1] , \y[0][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_3 \genblk1[1].element  ( 
        .clk(clk), .a({\a[7][7] , \a[7][6] , n147, \a[7][4] , \a[7][3] , 
        \a[7][2] , \a[7][1] , \a[7][0] , n105, \a[6][6] , n399, \a[6][4] , 
        n123, \a[6][2] , n148, \a[6][0] , n74, \a[5][6] , n139, \a[5][4] , n42, 
        \a[5][2] , n96, \a[5][0] , \a[4][7] , \a[4][6] , n397, \a[4][4] , n387, 
        \a[4][2] , \a[4][1] , \a[4][0] }), .x({n31, n93, n214, \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , n65, \x[2][6] , n215, 
        \x[2][4] , \x[2][3] , \x[2][2] , n87, \x[2][0] , n56, n27, \x[1][5] , 
        n6, \x[1][3] , \x[1][2] , n85, \x[1][0] , n44, n54, \x[0][5] , 
        \x[0][4] , n36, n67, n63, \x[0][0] }), .y({\y[1][15] , \y[1][14] , 
        \y[1][13] , \y[1][12] , \y[1][11] , \y[1][10] , \y[1][9] , \y[1][8] , 
        \y[1][7] , \y[1][6] , \y[1][5] , \y[1][4] , \y[1][3] , \y[1][2] , 
        \y[1][1] , \y[1][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_2 \genblk1[2].element  ( 
        .clk(clk), .a({\a[11][7] , \a[11][6] , n83, \a[11][4] , n403, 
        \a[11][2] , \a[11][1] , \a[11][0] , \a[10][7] , \a[10][6] , n76, 
        \a[10][4] , \a[10][3] , \a[10][2] , \a[10][1] , \a[10][0] , \a[9][7] , 
        \a[9][6] , \a[9][5] , \a[9][4] , \a[9][3] , \a[9][2] , \a[9][1] , 
        \a[9][0] , \a[8][7] , \a[8][6] , \a[8][5] , \a[8][4] , \a[8][3] , 
        \a[8][2] , \a[8][1] , \a[8][0] }), .x({n31, n93, n214, \x[3][4] , 
        \x[3][3] , \x[3][2] , n18, \x[3][0] , \x[2][7] , n29, n215, \x[2][4] , 
        \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , n56, \x[1][6] , \x[1][5] , 
        n6, n13, \x[1][2] , \x[1][1] , \x[1][0] , n44, n54, \x[0][5] , n25, 
        n36, n67, n63, \x[0][0] }), .y({\y[2][15] , \y[2][14] , \y[2][13] , 
        \y[2][12] , \y[2][11] , \y[2][10] , \y[2][9] , \y[2][8] , \y[2][7] , 
        \y[2][6] , \y[2][5] , \y[2][4] , \y[2][3] , \y[2][2] , \y[2][1] , 
        \y[2][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_1 \genblk1[3].element  ( 
        .clk(clk), .a({\a[15][7] , \a[15][6] , \a[15][5] , \a[15][4] , n395, 
        \a[15][2] , n141, \a[15][0] , \a[14][7] , \a[14][6] , \a[14][5] , 
        \a[14][4] , \a[14][3] , \a[14][2] , n401, \a[14][0] , n23, \a[13][6] , 
        \a[13][5] , \a[13][4] , \a[13][3] , \a[13][2] , \a[13][1] , \a[13][0] , 
        \a[12][7] , \a[12][6] , n391, \a[12][4] , n113, \a[12][2] , \a[12][1] , 
        \a[12][0] }), .x({\x[3][7] , n93, n214, \x[3][4] , \x[3][3] , 
        \x[3][2] , n18, \x[3][0] , n65, \x[2][6] , n215, \x[2][4] , \x[2][3] , 
        \x[2][2] , n87, \x[2][0] , \x[1][7] , n27, \x[1][5] , n6, \x[1][3] , 
        \x[1][2] , n85, \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , n25, n36, 
        n67, n63, \x[0][0] }), .y({\y[3][15] , \y[3][14] , \y[3][13] , 
        \y[3][12] , \y[3][11] , \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , 
        \y[3][6] , \y[3][5] , \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , 
        \y[3][0] }) );
  DFF_X2 \x_reg[1][2]  ( .D(n248), .CK(clk), .Q(\x[1][2] ) );
  DFF_X2 \x_reg[2][2]  ( .D(n240), .CK(clk), .Q(\x[2][2] ) );
  DFF_X2 \x_reg[3][2]  ( .D(n431), .CK(clk), .Q(\x[3][2] ) );
  DFF_X2 \x_reg[1][3]  ( .D(n247), .CK(clk), .Q(\x[1][3] ), .QN(n11) );
  DFF_X1 \a_reg[7][1]  ( .D(n329), .CK(clk), .Q(\a[7][1] ) );
  DFF_X2 \x_reg[3][3]  ( .D(n430), .CK(clk), .Q(\x[3][3] ) );
  DFF_X1 \a_reg[8][1]  ( .D(n321), .CK(clk), .Q(\a[8][1] ) );
  DFF_X1 \a_reg[13][3]  ( .D(n279), .CK(clk), .Q(\a[13][3] ) );
  DFF_X1 \a_reg[11][3]  ( .D(n295), .CK(clk), .Q(\a[11][3] ), .QN(n402) );
  DFF_X1 \a_reg[13][1]  ( .D(n281), .CK(clk), .Q(\a[13][1] ) );
  DFF_X1 \a_reg[14][1]  ( .D(n273), .CK(clk), .QN(n400) );
  DFF_X1 \a_reg[6][5]  ( .D(n333), .CK(clk), .Q(\a[6][5] ), .QN(n398) );
  DFF_X1 \a_reg[4][5]  ( .D(n349), .CK(clk), .Q(\a[4][5] ), .QN(n396) );
  DFF_X1 \a_reg[15][3]  ( .D(n263), .CK(clk), .Q(\a[15][3] ), .QN(n394) );
  DFF_X1 \a_reg[12][5]  ( .D(n285), .CK(clk), .Q(\a[12][5] ), .QN(n390) );
  DFF_X1 \a_reg[15][5]  ( .D(n261), .CK(clk), .Q(\a[15][5] ), .QN(n388) );
  DFF_X2 \x_reg[2][3]  ( .D(n239), .CK(clk), .Q(\x[2][3] ) );
  DFF_X1 \a_reg[14][3]  ( .D(n271), .CK(clk), .Q(\a[14][3] ) );
  DFF_X1 \a_reg[4][3]  ( .D(n351), .CK(clk), .QN(n230) );
  DFF_X1 \a_reg[13][5]  ( .D(n277), .CK(clk), .Q(\a[13][5] ) );
  DFF_X2 \x_reg[0][5]  ( .D(n253), .CK(clk), .Q(\x[0][5] ), .QN(n216) );
  DFF_X1 \a_reg[10][3]  ( .D(n303), .CK(clk), .Q(\a[10][3] ) );
  DFF_X1 \a_reg[1][5]  ( .D(n373), .CK(clk), .Q(\a[1][5] ), .QN(n7) );
  DFF_X1 \a_reg[0][3]  ( .D(n383), .CK(clk), .Q(\a[0][3] ) );
  DFF_X1 \a_reg[3][3]  ( .D(n359), .CK(clk), .Q(\a[3][3] ) );
  DFF_X1 \a_reg[7][3]  ( .D(n327), .CK(clk), .Q(\a[7][3] ), .QN(n33) );
  DFF_X1 \a_reg[3][5]  ( .D(n357), .CK(clk), .Q(\a[3][5] ) );
  DFF_X1 \a_reg[12][1]  ( .D(n289), .CK(clk), .Q(\a[12][1] ) );
  DFF_X1 \a_reg[14][5]  ( .D(n269), .CK(clk), .Q(\a[14][5] ) );
  DFF_X1 \a_reg[0][5]  ( .D(n381), .CK(clk), .Q(\a[0][5] ) );
  DFF_X2 \a_reg[15][7]  ( .D(n259), .CK(clk), .Q(\a[15][7] ) );
  DFF_X1 \a_reg[6][1]  ( .D(n337), .CK(clk), .Q(n148) );
  DFF_X1 \a_reg[7][5]  ( .D(n325), .CK(clk), .Q(\a[7][5] ), .QN(n142) );
  DFF_X2 \a_reg[2][7]  ( .D(n363), .CK(clk), .Q(\a[2][7] ) );
  DFF_X2 \a_reg[4][7]  ( .D(n347), .CK(clk), .Q(\a[4][7] ) );
  DFF_X1 \a_reg[15][1]  ( .D(n265), .CK(clk), .Q(\a[15][1] ), .QN(n140) );
  DFF_X2 \a_reg[4][1]  ( .D(n353), .CK(clk), .Q(\a[4][1] ), .QN(n404) );
  DFF_X1 \a_reg[5][5]  ( .D(n341), .CK(clk), .Q(\a[5][5] ), .QN(n138) );
  DFF_X1 \a_reg[2][5]  ( .D(n365), .CK(clk), .Q(\a[2][5] ), .QN(n132) );
  DFF_X1 \a_reg[0][7]  ( .D(n379), .CK(clk), .Q(\a[0][7] ) );
  DFF_X2 \x_reg[1][5]  ( .D(n245), .CK(clk), .Q(\x[1][5] ) );
  DFF_X1 \a_reg[1][7]  ( .D(n371), .CK(clk), .Q(\a[1][7] ), .QN(n124) );
  DFF_X1 \a_reg[0][1]  ( .D(n385), .CK(clk), .Q(\a[0][1] ) );
  DFF_X1 \a_reg[8][5]  ( .D(n317), .CK(clk), .Q(\a[8][5] ) );
  DFF_X2 \x_reg[3][4]  ( .D(n429), .CK(clk), .Q(\x[3][4] ) );
  DFF_X1 \a_reg[3][1]  ( .D(n361), .CK(clk), .Q(\a[3][1] ) );
  DFF_X2 \a_reg[8][7]  ( .D(n315), .CK(clk), .Q(\a[8][7] ) );
  DFF_X1 \a_reg[1][1]  ( .D(n377), .CK(clk), .Q(\a[1][1] ) );
  DFF_X1 \a_reg[6][3]  ( .D(n335), .CK(clk), .Q(\a[6][3] ), .QN(n122) );
  DFF_X1 \a_reg[3][7]  ( .D(n355), .CK(clk), .Q(\a[3][7] ), .QN(n114) );
  DFF_X2 \x_reg[2][4]  ( .D(n238), .CK(clk), .Q(\x[2][4] ) );
  DFF_X1 \a_reg[1][3]  ( .D(n375), .CK(clk), .Q(\a[1][3] ) );
  DFF_X1 \a_reg[12][3]  ( .D(n287), .CK(clk), .QN(n106) );
  DFF_X1 \a_reg[6][7]  ( .D(n331), .CK(clk), .Q(\a[6][7] ), .QN(n104) );
  DFF_X1 \a_reg[5][1]  ( .D(n345), .CK(clk), .Q(n96) );
  DFF_X1 \x_reg[3][6]  ( .D(n427), .CK(clk), .Q(\x[3][6] ), .QN(n92) );
  DFF_X1 \x_reg[2][1]  ( .D(n241), .CK(clk), .Q(\x[2][1] ), .QN(n86) );
  DFF_X1 \a_reg[8][3]  ( .D(n319), .CK(clk), .Q(\a[8][3] ), .QN(n392) );
  DFF_X1 \x_reg[1][1]  ( .D(n249), .CK(clk), .Q(\x[1][1] ), .QN(n84) );
  DFF_X1 \a_reg[11][5]  ( .D(n293), .CK(clk), .Q(\a[11][5] ), .QN(n77) );
  DFF_X1 \a_reg[10][5]  ( .D(n301), .CK(clk), .Q(\a[10][5] ), .QN(n75) );
  DFF_X1 \x_reg[0][2]  ( .D(n256), .CK(clk), .Q(\x[0][2] ), .QN(n66) );
  DFF_X1 \a_reg[9][5]  ( .D(n309), .CK(clk), .Q(\a[9][5] ) );
  DFF_X1 \x_reg[2][7]  ( .D(n235), .CK(clk), .Q(\x[2][7] ), .QN(n64) );
  DFF_X1 \a_reg[11][7]  ( .D(n291), .CK(clk), .Q(\a[11][7] ) );
  DFF_X1 \x_reg[0][1]  ( .D(n257), .CK(clk), .Q(\x[0][1] ), .QN(n57) );
  DFF_X1 \x_reg[1][7]  ( .D(n243), .CK(clk), .Q(\x[1][7] ), .QN(n55) );
  DFF_X1 \x_reg[0][6]  ( .D(n252), .CK(clk), .Q(\x[0][6] ), .QN(n53) );
  DFF_X1 \a_reg[5][3]  ( .D(n343), .CK(clk), .Q(\a[5][3] ), .QN(n37) );
  DFF_X1 \addr_y_reg[0]  ( .D(N101), .CK(clk), .Q(N24), .QN(n208) );
  DFF_X1 \a_reg[10][1]  ( .D(n305), .CK(clk), .Q(\a[10][1] ) );
  DFF_X1 \a_reg[2][2]  ( .D(n368), .CK(clk), .Q(\a[2][2] ) );
  DFF_X1 \a_reg[9][2]  ( .D(n312), .CK(clk), .Q(\a[9][2] ) );
  DFF_X1 \a_reg[4][4]  ( .D(n350), .CK(clk), .Q(\a[4][4] ) );
  DFF_X1 \a_reg[7][4]  ( .D(n326), .CK(clk), .Q(\a[7][4] ) );
  DFF_X1 \a_reg[14][2]  ( .D(n272), .CK(clk), .Q(\a[14][2] ) );
  DFF_X1 \a_reg[9][7]  ( .D(n307), .CK(clk), .Q(\a[9][7] ) );
  DFF_X1 \x_reg[2][6]  ( .D(n236), .CK(clk), .Q(\x[2][6] ), .QN(n28) );
  DFF_X1 \x_reg[1][6]  ( .D(n244), .CK(clk), .Q(\x[1][6] ), .QN(n26) );
  DFF_X1 \x_reg[0][4]  ( .D(n254), .CK(clk), .Q(\x[0][4] ), .QN(n24) );
  DFF_X2 \a_reg[14][7]  ( .D(n267), .CK(clk), .Q(\a[14][7] ) );
  DFF_X1 \a_reg[13][7]  ( .D(n275), .CK(clk), .Q(\a[13][7] ), .QN(n22) );
  DFF_X1 \x_reg[3][1]  ( .D(n432), .CK(clk), .Q(\x[3][1] ), .QN(n17) );
  DFF_X1 \x_reg[1][4]  ( .D(n246), .CK(clk), .Q(\x[1][4] ) );
  DFF_X1 \a_reg[2][3]  ( .D(n367), .CK(clk), .Q(\a[2][3] ) );
  DFF_X1 \a_reg[2][1]  ( .D(n369), .CK(clk), .Q(\a[2][1] ), .QN(n94) );
  DFF_X2 \a_reg[9][1]  ( .D(n313), .CK(clk), .Q(\a[9][1] ) );
  DFF_X2 \a_reg[9][3]  ( .D(n311), .CK(clk), .Q(\a[9][3] ) );
  DFF_X2 \a_reg[11][1]  ( .D(n297), .CK(clk), .Q(\a[11][1] ) );
  DFF_X1 \a_reg[11][0]  ( .D(n298), .CK(clk), .Q(\a[11][0] ) );
  DFF_X1 \a_reg[9][0]  ( .D(n314), .CK(clk), .Q(\a[9][0] ) );
  DFF_X1 \a_reg[7][6]  ( .D(n324), .CK(clk), .Q(\a[7][6] ) );
  INV_X2 U3 ( .A(n75), .ZN(n76) );
  AND2_X1 U4 ( .A1(N24), .A2(n3), .ZN(n1) );
  AND2_X1 U5 ( .A1(N25), .A2(n208), .ZN(n2) );
  AND2_X1 U6 ( .A1(n3), .A2(n208), .ZN(n4) );
  NOR3_X1 U7 ( .A1(n231), .A2(delay_timer[3]), .A3(n19), .ZN(n5) );
  BUF_X4 U8 ( .A(\x[1][4] ), .Z(n6) );
  INV_X1 U9 ( .A(n7), .ZN(n8) );
  INV_X1 U10 ( .A(n11), .ZN(n13) );
  CLKBUF_X1 U11 ( .A(n401), .Z(n14) );
  INV_X2 U12 ( .A(n17), .ZN(n18) );
  INV_X2 U13 ( .A(n22), .ZN(n23) );
  INV_X2 U14 ( .A(n24), .ZN(n25) );
  INV_X2 U15 ( .A(n26), .ZN(n27) );
  INV_X2 U16 ( .A(n28), .ZN(n29) );
  INV_X1 U17 ( .A(n30), .ZN(n31) );
  INV_X1 U18 ( .A(n33), .ZN(n34) );
  INV_X2 U19 ( .A(n35), .ZN(n36) );
  INV_X2 U20 ( .A(n37), .ZN(n42) );
  INV_X2 U21 ( .A(n43), .ZN(n44) );
  INV_X1 U22 ( .A(n45), .ZN(n46) );
  INV_X2 U23 ( .A(n53), .ZN(n54) );
  INV_X2 U24 ( .A(n55), .ZN(n56) );
  INV_X2 U25 ( .A(n57), .ZN(n63) );
  INV_X2 U26 ( .A(n64), .ZN(n65) );
  INV_X2 U27 ( .A(n66), .ZN(n67) );
  INV_X2 U28 ( .A(n73), .ZN(n74) );
  INV_X2 U29 ( .A(n77), .ZN(n83) );
  INV_X2 U30 ( .A(n84), .ZN(n85) );
  INV_X2 U31 ( .A(n86), .ZN(n87) );
  INV_X2 U32 ( .A(n92), .ZN(n93) );
  INV_X1 U33 ( .A(n94), .ZN(n95) );
  INV_X2 U34 ( .A(n104), .ZN(n105) );
  INV_X2 U35 ( .A(n106), .ZN(n113) );
  INV_X2 U36 ( .A(n114), .ZN(n115) );
  INV_X2 U37 ( .A(n122), .ZN(n123) );
  INV_X2 U38 ( .A(n124), .ZN(n131) );
  INV_X2 U39 ( .A(n132), .ZN(n133) );
  INV_X2 U40 ( .A(n138), .ZN(n139) );
  INV_X2 U41 ( .A(n140), .ZN(n141) );
  INV_X2 U42 ( .A(n142), .ZN(n147) );
  INV_X1 U43 ( .A(data_in[6]), .ZN(n440) );
  INV_X1 U44 ( .A(data_in[7]), .ZN(n439) );
  INV_X1 U45 ( .A(n208), .ZN(n213) );
  OAI21_X1 U46 ( .B1(n443), .B2(n125), .A(n130), .ZN(n255) );
  OAI21_X1 U47 ( .B1(n439), .B2(n125), .A(n126), .ZN(n251) );
  OAI21_X1 U48 ( .B1(n441), .B2(n125), .A(n128), .ZN(n253) );
  NAND2_X1 U49 ( .A1(n217), .A2(n125), .ZN(n128) );
  OAI21_X1 U50 ( .B1(n441), .B2(n107), .A(n110), .ZN(n237) );
  NAND2_X1 U51 ( .A1(n215), .A2(n107), .ZN(n110) );
  INV_X1 U52 ( .A(n227), .ZN(n435) );
  OAI21_X1 U53 ( .B1(n78), .B2(n47), .A(n436), .ZN(n227) );
  NAND3_X1 U54 ( .A1(addr_x[0]), .A2(n15), .A3(en_x), .ZN(n116) );
  NOR4_X1 U55 ( .A1(delay_timer[3]), .A2(delay_timer[2]), .A3(delay_timer[1]), 
        .A4(n21), .ZN(of_delay) );
  NAND3_X1 U56 ( .A1(n15), .A2(n16), .A3(en_x), .ZN(n125) );
  NAND3_X1 U57 ( .A1(addr_x[1]), .A2(n16), .A3(en_x), .ZN(n107) );
  NOR3_X1 U58 ( .A1(n225), .A2(n10), .A3(n9), .ZN(N114) );
  NOR2_X1 U59 ( .A1(n12), .A2(addr_a[0]), .ZN(n78) );
  NOR2_X1 U60 ( .A1(n15), .A2(n16), .ZN(N115) );
  AOI21_X1 U61 ( .B1(n20), .B2(n438), .A(N108), .ZN(n232) );
  AOI21_X1 U62 ( .B1(n436), .B2(n12), .A(N89), .ZN(n222) );
  OAI21_X1 U63 ( .B1(n442), .B2(n125), .A(n129), .ZN(n254) );
  NAND2_X1 U64 ( .A1(n25), .A2(n125), .ZN(n129) );
  OAI21_X1 U65 ( .B1(n442), .B2(n107), .A(n111), .ZN(n238) );
  NAND2_X1 U66 ( .A1(\x[2][4] ), .A2(n107), .ZN(n111) );
  NOR2_X1 U67 ( .A1(addr_a[0]), .A2(addr_a[1]), .ZN(n58) );
  OAI22_X1 U68 ( .A1(n232), .A2(n19), .B1(delay_timer[2]), .B2(n231), .ZN(N110) );
  NOR2_X1 U69 ( .A1(clr_addr_y), .A2(n234), .ZN(N102) );
  XNOR2_X1 U70 ( .A(N25), .B(N24), .ZN(n234) );
  OAI22_X1 U71 ( .A1(n222), .A2(n9), .B1(clr_addr_a), .B2(n223), .ZN(N92) );
  AOI22_X1 U72 ( .A1(n224), .A2(n425), .B1(addr_a[3]), .B2(n10), .ZN(n223) );
  NOR2_X1 U73 ( .A1(addr_a[3]), .A2(n10), .ZN(n224) );
  OAI22_X1 U74 ( .A1(n222), .A2(n10), .B1(n225), .B2(n226), .ZN(N91) );
  NAND2_X1 U75 ( .A1(n10), .A2(n436), .ZN(n226) );
  OAI21_X1 U76 ( .B1(n439), .B2(n162), .A(n163), .ZN(n283) );
  NAND2_X1 U77 ( .A1(\a[12][7] ), .A2(n162), .ZN(n163) );
  OAI21_X1 U78 ( .B1(n439), .B2(n200), .A(n201), .ZN(n315) );
  NAND2_X1 U79 ( .A1(\a[8][7] ), .A2(n200), .ZN(n201) );
  OAI21_X1 U80 ( .B1(n439), .B2(n191), .A(n192), .ZN(n307) );
  NAND2_X1 U81 ( .A1(n29), .A2(n107), .ZN(n109) );
  INV_X1 U82 ( .A(n216), .ZN(n217) );
  NOR2_X1 U83 ( .A1(clr_delay), .A2(delay_timer[0]), .ZN(N108) );
  NOR2_X1 U84 ( .A1(addr_a[0]), .A2(clr_addr_a), .ZN(N89) );
  OAI21_X1 U85 ( .B1(n38), .B2(n439), .A(n39), .ZN(n339) );
  NAND2_X1 U86 ( .A1(\a[5][7] ), .A2(n38), .ZN(n39) );
  OAI21_X1 U87 ( .B1(n38), .B2(n441), .A(n41), .ZN(n341) );
  OAI21_X1 U88 ( .B1(n441), .B2(n69), .A(n72), .ZN(n365) );
  OAI21_X1 U89 ( .B1(n441), .B2(n88), .A(n91), .ZN(n381) );
  OAI21_X1 U90 ( .B1(n442), .B2(n116), .A(n120), .ZN(n246) );
  NAND2_X1 U91 ( .A1(n6), .A2(n116), .ZN(n120) );
  OAI21_X1 U92 ( .B1(n441), .B2(n116), .A(n119), .ZN(n245) );
  NAND2_X1 U93 ( .A1(\x[1][5] ), .A2(n116), .ZN(n119) );
  OAI21_X1 U94 ( .B1(n440), .B2(n116), .A(n118), .ZN(n244) );
  NAND2_X1 U95 ( .A1(n27), .A2(n116), .ZN(n118) );
  OAI21_X1 U96 ( .B1(n443), .B2(n116), .A(n121), .ZN(n247) );
  NAND2_X1 U97 ( .A1(n13), .A2(n116), .ZN(n121) );
  OAI21_X1 U98 ( .B1(n439), .B2(n116), .A(n117), .ZN(n243) );
  NAND2_X1 U99 ( .A1(n56), .A2(n116), .ZN(n117) );
  OAI21_X1 U100 ( .B1(n32), .B2(n440), .A(n219), .ZN(n332) );
  NAND2_X1 U101 ( .A1(\a[6][6] ), .A2(n32), .ZN(n219) );
  OAI21_X1 U102 ( .B1(n32), .B2(n439), .A(n218), .ZN(n331) );
  OAI21_X1 U103 ( .B1(n440), .B2(n125), .A(n127), .ZN(n252) );
  AND2_X1 U104 ( .A1(addr_a[0]), .A2(n12), .ZN(n47) );
  OAI21_X1 U105 ( .B1(n439), .B2(n107), .A(n108), .ZN(n235) );
  OAI21_X1 U106 ( .B1(n440), .B2(n69), .A(n71), .ZN(n364) );
  NAND2_X1 U107 ( .A1(\a[2][6] ), .A2(n69), .ZN(n71) );
  OAI21_X1 U108 ( .B1(n439), .B2(n69), .A(n70), .ZN(n363) );
  OAI21_X1 U109 ( .B1(n439), .B2(n88), .A(n89), .ZN(n379) );
  OAI21_X1 U110 ( .B1(n440), .B2(n182), .A(n184), .ZN(n300) );
  NAND2_X1 U111 ( .A1(\a[10][6] ), .A2(n182), .ZN(n184) );
  OAI21_X1 U112 ( .B1(n439), .B2(n182), .A(n183), .ZN(n299) );
  NAND2_X1 U113 ( .A1(n46), .A2(n182), .ZN(n183) );
  OAI21_X1 U114 ( .B1(n440), .B2(n172), .A(n174), .ZN(n292) );
  NAND2_X1 U115 ( .A1(\a[11][6] ), .A2(n172), .ZN(n174) );
  NAND2_X1 U116 ( .A1(addr_a[0]), .A2(addr_a[1]), .ZN(n225) );
  OAI21_X1 U117 ( .B1(n439), .B2(n134), .A(n135), .ZN(n259) );
  OAI21_X1 U118 ( .B1(n439), .B2(n143), .A(n144), .ZN(n267) );
  OAI21_X1 U119 ( .B1(n439), .B2(n49), .A(n50), .ZN(n347) );
  OAI21_X1 U120 ( .B1(n440), .B2(n209), .A(n211), .ZN(n324) );
  NAND2_X1 U121 ( .A1(\a[7][6] ), .A2(n209), .ZN(n211) );
  OAI21_X1 U122 ( .B1(n439), .B2(n209), .A(n210), .ZN(n323) );
  OAI21_X1 U123 ( .B1(n440), .B2(n59), .A(n61), .ZN(n356) );
  NAND2_X1 U124 ( .A1(\a[3][6] ), .A2(n59), .ZN(n61) );
  OAI21_X1 U125 ( .B1(n439), .B2(n59), .A(n60), .ZN(n355) );
  OAI21_X1 U126 ( .B1(n440), .B2(n79), .A(n81), .ZN(n372) );
  NAND2_X1 U127 ( .A1(\a[1][6] ), .A2(n79), .ZN(n81) );
  OAI21_X1 U128 ( .B1(n439), .B2(n79), .A(n80), .ZN(n371) );
  OAI21_X1 U129 ( .B1(n440), .B2(n191), .A(n193), .ZN(n308) );
  NAND2_X1 U130 ( .A1(\a[9][6] ), .A2(n191), .ZN(n193) );
  OAI21_X1 U131 ( .B1(n440), .B2(n153), .A(n155), .ZN(n276) );
  NAND2_X1 U132 ( .A1(\a[13][6] ), .A2(n153), .ZN(n155) );
  OAI21_X1 U133 ( .B1(n440), .B2(n88), .A(n90), .ZN(n380) );
  NAND2_X1 U134 ( .A1(\a[0][6] ), .A2(n88), .ZN(n90) );
  OAI21_X1 U135 ( .B1(n440), .B2(n162), .A(n164), .ZN(n284) );
  NAND2_X1 U136 ( .A1(\a[12][6] ), .A2(n162), .ZN(n164) );
  OAI21_X1 U137 ( .B1(n440), .B2(n200), .A(n202), .ZN(n316) );
  NAND2_X1 U138 ( .A1(\a[8][6] ), .A2(n200), .ZN(n202) );
  OAI21_X1 U139 ( .B1(n439), .B2(n172), .A(n173), .ZN(n291) );
  NAND2_X1 U140 ( .A1(\a[11][7] ), .A2(n172), .ZN(n173) );
  OAI21_X1 U141 ( .B1(n38), .B2(n440), .A(n40), .ZN(n340) );
  NAND2_X1 U142 ( .A1(\a[5][6] ), .A2(n38), .ZN(n40) );
  INV_X1 U143 ( .A(clr_addr_a), .ZN(n436) );
  OAI21_X1 U144 ( .B1(n440), .B2(n134), .A(n136), .ZN(n260) );
  NAND2_X1 U145 ( .A1(\a[15][6] ), .A2(n134), .ZN(n136) );
  OAI21_X1 U146 ( .B1(n440), .B2(n143), .A(n145), .ZN(n268) );
  NAND2_X1 U147 ( .A1(\a[14][6] ), .A2(n143), .ZN(n145) );
  OAI21_X1 U148 ( .B1(n440), .B2(n49), .A(n51), .ZN(n348) );
  NAND2_X1 U149 ( .A1(\a[4][6] ), .A2(n49), .ZN(n51) );
  AND2_X1 U150 ( .A1(n97), .A2(n10), .ZN(n68) );
  AND2_X1 U151 ( .A1(n171), .A2(n10), .ZN(n181) );
  AND2_X1 U152 ( .A1(N24), .A2(N25), .ZN(N116) );
  AND2_X1 U153 ( .A1(addr_a[2]), .A2(n97), .ZN(n48) );
  NOR2_X1 U154 ( .A1(clr_delay), .A2(n233), .ZN(N109) );
  XNOR2_X1 U155 ( .A(delay_timer[0]), .B(delay_timer[1]), .ZN(n233) );
  INV_X1 U156 ( .A(clr_delay), .ZN(n438) );
  NOR2_X1 U157 ( .A1(clr_addr_y), .A2(N24), .ZN(N101) );
  NOR2_X1 U158 ( .A1(clr_addr_x), .A2(n221), .ZN(N97) );
  XNOR2_X1 U159 ( .A(addr_x[1]), .B(addr_x[0]), .ZN(n221) );
  NOR2_X1 U160 ( .A1(clr_addr_x), .A2(addr_x[0]), .ZN(N96) );
  AND2_X1 U161 ( .A1(n171), .A2(addr_a[2]), .ZN(n152) );
  AND2_X1 U162 ( .A1(en_a), .A2(n9), .ZN(n97) );
  AND2_X1 U163 ( .A1(addr_a[3]), .A2(en_a), .ZN(n171) );
  INV_X1 U164 ( .A(n102), .ZN(n429) );
  AOI22_X1 U165 ( .A1(data_in[4]), .A2(n434), .B1(n99), .B2(\x[3][4] ), .ZN(
        n102) );
  INV_X1 U166 ( .A(n100), .ZN(n427) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n434), .B1(n99), .B2(n93), .ZN(n100) );
  INV_X1 U168 ( .A(n98), .ZN(n426) );
  INV_X1 U169 ( .A(n101), .ZN(n428) );
  AOI22_X1 U170 ( .A1(data_in[5]), .A2(n434), .B1(n99), .B2(n214), .ZN(n101)
         );
  INV_X1 U171 ( .A(n103), .ZN(n430) );
  AOI22_X1 U172 ( .A1(data_in[3]), .A2(n434), .B1(n99), .B2(\x[3][3] ), .ZN(
        n103) );
  INV_X1 U173 ( .A(n228), .ZN(n437) );
  AOI21_X1 U174 ( .B1(n229), .B2(delay_timer[3]), .A(n5), .ZN(n228) );
  OAI21_X1 U175 ( .B1(clr_delay), .B2(delay_timer[2]), .A(n232), .ZN(n229) );
  INV_X1 U176 ( .A(data_in[5]), .ZN(n441) );
  MUX2_X1 U177 ( .A(\y[2][0] ), .B(\y[3][0] ), .S(n213), .Z(n149) );
  MUX2_X1 U178 ( .A(\y[0][0] ), .B(\y[1][0] ), .S(n213), .Z(n150) );
  MUX2_X1 U179 ( .A(n150), .B(n149), .S(N25), .Z(N83) );
  MUX2_X1 U180 ( .A(\y[2][1] ), .B(\y[3][1] ), .S(n213), .Z(n151) );
  MUX2_X1 U181 ( .A(\y[0][1] ), .B(\y[1][1] ), .S(n213), .Z(n157) );
  MUX2_X1 U182 ( .A(n157), .B(n151), .S(N25), .Z(N82) );
  MUX2_X1 U183 ( .A(\y[2][2] ), .B(\y[3][2] ), .S(n213), .Z(n158) );
  MUX2_X1 U184 ( .A(\y[0][2] ), .B(\y[1][2] ), .S(n213), .Z(n159) );
  MUX2_X1 U185 ( .A(n159), .B(n158), .S(N25), .Z(N81) );
  MUX2_X1 U186 ( .A(\y[2][3] ), .B(\y[3][3] ), .S(n213), .Z(n160) );
  MUX2_X1 U187 ( .A(\y[0][3] ), .B(\y[1][3] ), .S(n213), .Z(n161) );
  MUX2_X1 U188 ( .A(n161), .B(n160), .S(N25), .Z(N80) );
  MUX2_X1 U189 ( .A(\y[2][4] ), .B(\y[3][4] ), .S(n213), .Z(n166) );
  MUX2_X1 U190 ( .A(\y[0][4] ), .B(\y[1][4] ), .S(n213), .Z(n167) );
  MUX2_X1 U191 ( .A(n167), .B(n166), .S(N25), .Z(N79) );
  MUX2_X1 U192 ( .A(\y[2][5] ), .B(\y[3][5] ), .S(n213), .Z(n168) );
  MUX2_X1 U193 ( .A(\y[0][5] ), .B(\y[1][5] ), .S(n213), .Z(n169) );
  MUX2_X1 U194 ( .A(n169), .B(n168), .S(N25), .Z(N78) );
  MUX2_X1 U195 ( .A(\y[2][6] ), .B(\y[3][6] ), .S(n213), .Z(n170) );
  MUX2_X1 U196 ( .A(\y[0][6] ), .B(\y[1][6] ), .S(n213), .Z(n176) );
  MUX2_X1 U197 ( .A(n176), .B(n170), .S(N25), .Z(N77) );
  MUX2_X1 U198 ( .A(\y[2][7] ), .B(\y[3][7] ), .S(N24), .Z(n177) );
  MUX2_X1 U199 ( .A(\y[0][7] ), .B(\y[1][7] ), .S(N24), .Z(n178) );
  MUX2_X1 U200 ( .A(n178), .B(n177), .S(N25), .Z(N76) );
  MUX2_X1 U201 ( .A(\y[2][8] ), .B(\y[3][8] ), .S(n213), .Z(n179) );
  MUX2_X1 U202 ( .A(\y[0][8] ), .B(\y[1][8] ), .S(N24), .Z(n180) );
  MUX2_X1 U203 ( .A(n180), .B(n179), .S(N25), .Z(N75) );
  MUX2_X1 U204 ( .A(\y[2][9] ), .B(\y[3][9] ), .S(N24), .Z(n186) );
  MUX2_X1 U205 ( .A(\y[0][9] ), .B(\y[1][9] ), .S(n213), .Z(n187) );
  MUX2_X1 U206 ( .A(n187), .B(n186), .S(N25), .Z(N74) );
  MUX2_X1 U207 ( .A(\y[2][10] ), .B(\y[3][10] ), .S(n213), .Z(n188) );
  MUX2_X1 U208 ( .A(\y[0][10] ), .B(\y[1][10] ), .S(N24), .Z(n189) );
  MUX2_X1 U209 ( .A(n189), .B(n188), .S(N25), .Z(N73) );
  MUX2_X1 U210 ( .A(\y[2][11] ), .B(\y[3][11] ), .S(n213), .Z(n190) );
  MUX2_X1 U211 ( .A(\y[0][11] ), .B(\y[1][11] ), .S(N24), .Z(n195) );
  MUX2_X1 U212 ( .A(n195), .B(n190), .S(N25), .Z(N72) );
  NAND2_X1 U213 ( .A1(n196), .A2(n197), .ZN(N71) );
  AOI22_X1 U214 ( .A1(\y[1][12] ), .A2(n1), .B1(\y[3][12] ), .B2(N116), .ZN(
        n197) );
  AOI22_X1 U215 ( .A1(\y[0][12] ), .A2(n4), .B1(\y[2][12] ), .B2(n2), .ZN(n196) );
  NAND2_X1 U216 ( .A1(n198), .A2(n199), .ZN(N70) );
  AOI22_X1 U217 ( .A1(\y[1][13] ), .A2(n1), .B1(\y[3][13] ), .B2(N116), .ZN(
        n199) );
  AOI22_X1 U218 ( .A1(\y[0][13] ), .A2(n4), .B1(\y[2][13] ), .B2(n2), .ZN(n198) );
  NAND2_X1 U219 ( .A1(n205), .A2(n204), .ZN(N69) );
  AOI22_X1 U220 ( .A1(\y[1][14] ), .A2(n1), .B1(\y[3][14] ), .B2(N116), .ZN(
        n205) );
  AOI22_X1 U221 ( .A1(\y[0][14] ), .A2(n4), .B1(\y[2][14] ), .B2(n2), .ZN(n204) );
  NAND2_X1 U222 ( .A1(n207), .A2(n206), .ZN(N68) );
  AOI22_X1 U223 ( .A1(\y[1][15] ), .A2(n1), .B1(\y[3][15] ), .B2(N116), .ZN(
        n207) );
  AOI22_X1 U224 ( .A1(\y[0][15] ), .A2(n4), .B1(\y[2][15] ), .B2(n2), .ZN(n206) );
  BUF_X4 U225 ( .A(\x[3][5] ), .Z(n214) );
  OAI21_X1 U226 ( .B1(n439), .B2(n153), .A(n154), .ZN(n275) );
  OAI21_X1 U227 ( .B1(n441), .B2(n59), .A(n62), .ZN(n357) );
  INV_X1 U228 ( .A(n388), .ZN(n389) );
  INV_X1 U229 ( .A(n398), .ZN(n399) );
  NAND2_X1 U230 ( .A1(\a[4][7] ), .A2(n49), .ZN(n50) );
  NAND2_X1 U231 ( .A1(\a[14][7] ), .A2(n143), .ZN(n144) );
  NAND2_X1 U232 ( .A1(\a[0][7] ), .A2(n88), .ZN(n89) );
  OAI21_X1 U233 ( .B1(n441), .B2(n79), .A(n82), .ZN(n373) );
  NAND2_X1 U234 ( .A1(\a[3][7] ), .A2(n59), .ZN(n60) );
  NAND2_X1 U235 ( .A1(\a[6][7] ), .A2(n32), .ZN(n218) );
  NAND2_X1 U236 ( .A1(\a[2][7] ), .A2(n69), .ZN(n70) );
  NAND2_X1 U237 ( .A1(\a[9][7] ), .A2(n191), .ZN(n192) );
  BUF_X4 U238 ( .A(\x[2][5] ), .Z(n215) );
  OAI21_X1 U239 ( .B1(n32), .B2(n441), .A(n220), .ZN(n333) );
  NAND2_X1 U240 ( .A1(\a[1][7] ), .A2(n79), .ZN(n80) );
  INV_X2 U241 ( .A(n230), .ZN(n387) );
  OAI21_X1 U242 ( .B1(n441), .B2(n143), .A(n146), .ZN(n269) );
  OAI21_X1 U243 ( .B1(n443), .B2(n107), .A(n112), .ZN(n239) );
  NAND2_X1 U244 ( .A1(n54), .A2(n125), .ZN(n127) );
  OAI21_X1 U245 ( .B1(n440), .B2(n107), .A(n109), .ZN(n236) );
  OAI21_X1 U246 ( .B1(n441), .B2(n153), .A(n156), .ZN(n277) );
  OAI21_X1 U247 ( .B1(n441), .B2(n209), .A(n212), .ZN(n325) );
  OAI21_X1 U248 ( .B1(n441), .B2(n182), .A(n185), .ZN(n301) );
  INV_X2 U249 ( .A(n390), .ZN(n391) );
  OAI21_X1 U250 ( .B1(n441), .B2(n162), .A(n165), .ZN(n285) );
  INV_X1 U251 ( .A(n392), .ZN(n393) );
  INV_X2 U252 ( .A(n394), .ZN(n395) );
  INV_X2 U253 ( .A(n396), .ZN(n397) );
  OAI21_X1 U254 ( .B1(n441), .B2(n49), .A(n52), .ZN(n349) );
  OAI21_X1 U255 ( .B1(n441), .B2(n134), .A(n137), .ZN(n261) );
  OAI21_X1 U256 ( .B1(n441), .B2(n200), .A(n203), .ZN(n317) );
  INV_X2 U257 ( .A(n400), .ZN(n401) );
  NAND2_X1 U258 ( .A1(\a[7][7] ), .A2(n209), .ZN(n210) );
  INV_X2 U259 ( .A(n402), .ZN(n403) );
  NAND2_X1 U260 ( .A1(\a[15][7] ), .A2(n134), .ZN(n135) );
  OAI21_X1 U261 ( .B1(n441), .B2(n191), .A(n194), .ZN(n309) );
  NAND2_X1 U262 ( .A1(n44), .A2(n125), .ZN(n126) );
  NAND2_X1 U263 ( .A1(\a[13][7] ), .A2(n153), .ZN(n154) );
  NAND2_X1 U264 ( .A1(\a[4][5] ), .A2(n49), .ZN(n52) );
  OAI21_X1 U265 ( .B1(n441), .B2(n172), .A(n175), .ZN(n293) );
  NAND2_X1 U266 ( .A1(\a[14][5] ), .A2(n143), .ZN(n146) );
  NAND2_X1 U267 ( .A1(\x[2][3] ), .A2(n107), .ZN(n112) );
  INV_X1 U268 ( .A(n404), .ZN(n405) );
  NAND2_X1 U269 ( .A1(\a[12][5] ), .A2(n162), .ZN(n165) );
  AOI22_X1 U270 ( .A1(data_in[7]), .A2(n434), .B1(n99), .B2(\x[3][7] ), .ZN(
        n98) );
  NAND2_X1 U271 ( .A1(n65), .A2(n107), .ZN(n108) );
  NAND2_X1 U272 ( .A1(\a[8][5] ), .A2(n200), .ZN(n203) );
  NAND2_X1 U273 ( .A1(\a[10][5] ), .A2(n182), .ZN(n185) );
  NAND2_X1 U274 ( .A1(n36), .A2(n125), .ZN(n130) );
  NAND2_X1 U275 ( .A1(\a[0][5] ), .A2(n88), .ZN(n91) );
  NAND2_X1 U276 ( .A1(\a[2][5] ), .A2(n69), .ZN(n72) );
  NAND2_X1 U277 ( .A1(\a[6][5] ), .A2(n32), .ZN(n220) );
  NAND2_X1 U278 ( .A1(\a[9][5] ), .A2(n191), .ZN(n194) );
  NAND2_X1 U279 ( .A1(\a[5][5] ), .A2(n38), .ZN(n41) );
  NAND2_X1 U280 ( .A1(\a[7][5] ), .A2(n209), .ZN(n212) );
  NAND2_X1 U281 ( .A1(n8), .A2(n79), .ZN(n82) );
  NAND2_X1 U282 ( .A1(\a[13][5] ), .A2(n153), .ZN(n156) );
  NAND2_X1 U283 ( .A1(\a[3][5] ), .A2(n59), .ZN(n62) );
  NAND2_X1 U284 ( .A1(n389), .A2(n134), .ZN(n137) );
  NAND2_X1 U285 ( .A1(\a[11][5] ), .A2(n172), .ZN(n175) );
  NAND2_X1 U286 ( .A1(en_a), .A2(N114), .ZN(n134) );
  INV_X1 U287 ( .A(n134), .ZN(n406) );
  MUX2_X1 U288 ( .A(\a[15][4] ), .B(data_in[4]), .S(n406), .Z(n262) );
  MUX2_X1 U289 ( .A(\a[15][3] ), .B(data_in[3]), .S(n406), .Z(n263) );
  MUX2_X1 U290 ( .A(\a[15][2] ), .B(data_in[2]), .S(n406), .Z(n264) );
  MUX2_X1 U291 ( .A(\a[15][1] ), .B(data_in[1]), .S(n406), .Z(n265) );
  MUX2_X1 U292 ( .A(\a[15][0] ), .B(data_in[0]), .S(n406), .Z(n266) );
  NAND2_X1 U293 ( .A1(n152), .A2(n78), .ZN(n143) );
  INV_X1 U294 ( .A(n143), .ZN(n407) );
  MUX2_X1 U295 ( .A(\a[14][4] ), .B(data_in[4]), .S(n407), .Z(n270) );
  MUX2_X1 U296 ( .A(\a[14][3] ), .B(data_in[3]), .S(n407), .Z(n271) );
  MUX2_X1 U297 ( .A(\a[14][2] ), .B(data_in[2]), .S(n407), .Z(n272) );
  MUX2_X1 U298 ( .A(n14), .B(data_in[1]), .S(n407), .Z(n273) );
  MUX2_X1 U299 ( .A(\a[14][0] ), .B(data_in[0]), .S(n407), .Z(n274) );
  NAND2_X1 U300 ( .A1(n152), .A2(n47), .ZN(n153) );
  INV_X1 U301 ( .A(n153), .ZN(n408) );
  MUX2_X1 U302 ( .A(\a[13][4] ), .B(data_in[4]), .S(n408), .Z(n278) );
  MUX2_X1 U303 ( .A(\a[13][3] ), .B(data_in[3]), .S(n408), .Z(n279) );
  MUX2_X1 U304 ( .A(\a[13][2] ), .B(data_in[2]), .S(n408), .Z(n280) );
  MUX2_X1 U305 ( .A(\a[13][1] ), .B(data_in[1]), .S(n408), .Z(n281) );
  MUX2_X1 U306 ( .A(\a[13][0] ), .B(data_in[0]), .S(n408), .Z(n282) );
  NAND2_X1 U307 ( .A1(n152), .A2(n58), .ZN(n162) );
  INV_X1 U308 ( .A(n162), .ZN(n409) );
  MUX2_X1 U309 ( .A(\a[12][4] ), .B(data_in[4]), .S(n409), .Z(n286) );
  MUX2_X1 U310 ( .A(n113), .B(data_in[3]), .S(n409), .Z(n287) );
  MUX2_X1 U311 ( .A(\a[12][2] ), .B(data_in[2]), .S(n409), .Z(n288) );
  MUX2_X1 U312 ( .A(\a[12][1] ), .B(data_in[1]), .S(n409), .Z(n289) );
  MUX2_X1 U313 ( .A(\a[12][0] ), .B(data_in[0]), .S(n409), .Z(n290) );
  NAND2_X1 U314 ( .A1(en_x), .A2(N115), .ZN(n99) );
  INV_X1 U315 ( .A(n99), .ZN(n434) );
  MUX2_X1 U316 ( .A(\x[3][2] ), .B(data_in[2]), .S(n434), .Z(n431) );
  MUX2_X1 U317 ( .A(n18), .B(data_in[1]), .S(n434), .Z(n432) );
  MUX2_X1 U318 ( .A(\x[3][0] ), .B(data_in[0]), .S(n434), .Z(n433) );
  INV_X1 U319 ( .A(n107), .ZN(n410) );
  MUX2_X1 U320 ( .A(\x[2][2] ), .B(data_in[2]), .S(n410), .Z(n240) );
  MUX2_X1 U321 ( .A(n87), .B(data_in[1]), .S(n410), .Z(n241) );
  MUX2_X1 U322 ( .A(\x[2][0] ), .B(data_in[0]), .S(n410), .Z(n242) );
  INV_X1 U323 ( .A(n116), .ZN(n411) );
  MUX2_X1 U324 ( .A(\x[1][2] ), .B(data_in[2]), .S(n411), .Z(n248) );
  MUX2_X1 U325 ( .A(n85), .B(data_in[1]), .S(n411), .Z(n249) );
  MUX2_X1 U326 ( .A(\x[1][0] ), .B(data_in[0]), .S(n411), .Z(n250) );
  INV_X1 U327 ( .A(n125), .ZN(n412) );
  MUX2_X1 U328 ( .A(n67), .B(data_in[2]), .S(n412), .Z(n256) );
  MUX2_X1 U329 ( .A(n63), .B(data_in[1]), .S(n412), .Z(n257) );
  MUX2_X1 U330 ( .A(\x[0][0] ), .B(data_in[0]), .S(n412), .Z(n258) );
  INV_X1 U331 ( .A(n225), .ZN(n425) );
  NAND2_X1 U332 ( .A1(n181), .A2(n425), .ZN(n172) );
  INV_X1 U333 ( .A(n172), .ZN(n413) );
  MUX2_X1 U334 ( .A(\a[11][4] ), .B(data_in[4]), .S(n413), .Z(n294) );
  MUX2_X1 U335 ( .A(\a[11][3] ), .B(data_in[3]), .S(n413), .Z(n295) );
  MUX2_X1 U336 ( .A(\a[11][2] ), .B(data_in[2]), .S(n413), .Z(n296) );
  MUX2_X1 U337 ( .A(\a[11][1] ), .B(data_in[1]), .S(n413), .Z(n297) );
  MUX2_X1 U338 ( .A(\a[11][0] ), .B(data_in[0]), .S(n413), .Z(n298) );
  NAND2_X1 U339 ( .A1(n181), .A2(n78), .ZN(n182) );
  INV_X1 U340 ( .A(n182), .ZN(n414) );
  MUX2_X1 U341 ( .A(\a[10][4] ), .B(data_in[4]), .S(n414), .Z(n302) );
  MUX2_X1 U342 ( .A(\a[10][3] ), .B(data_in[3]), .S(n414), .Z(n303) );
  MUX2_X1 U343 ( .A(\a[10][2] ), .B(data_in[2]), .S(n414), .Z(n304) );
  MUX2_X1 U344 ( .A(\a[10][1] ), .B(data_in[1]), .S(n414), .Z(n305) );
  MUX2_X1 U345 ( .A(\a[10][0] ), .B(data_in[0]), .S(n414), .Z(n306) );
  NAND2_X1 U346 ( .A1(n181), .A2(n47), .ZN(n191) );
  INV_X1 U347 ( .A(n191), .ZN(n415) );
  MUX2_X1 U348 ( .A(\a[9][4] ), .B(data_in[4]), .S(n415), .Z(n310) );
  MUX2_X1 U349 ( .A(\a[9][3] ), .B(data_in[3]), .S(n415), .Z(n311) );
  MUX2_X1 U350 ( .A(\a[9][2] ), .B(data_in[2]), .S(n415), .Z(n312) );
  MUX2_X1 U351 ( .A(\a[9][1] ), .B(data_in[1]), .S(n415), .Z(n313) );
  MUX2_X1 U352 ( .A(\a[9][0] ), .B(data_in[0]), .S(n415), .Z(n314) );
  NAND2_X1 U353 ( .A1(n181), .A2(n58), .ZN(n200) );
  INV_X1 U354 ( .A(n200), .ZN(n416) );
  MUX2_X1 U355 ( .A(\a[8][4] ), .B(data_in[4]), .S(n416), .Z(n318) );
  MUX2_X1 U356 ( .A(n393), .B(data_in[3]), .S(n416), .Z(n319) );
  MUX2_X1 U357 ( .A(\a[8][2] ), .B(data_in[2]), .S(n416), .Z(n320) );
  MUX2_X1 U358 ( .A(\a[8][1] ), .B(data_in[1]), .S(n416), .Z(n321) );
  MUX2_X1 U359 ( .A(\a[8][0] ), .B(data_in[0]), .S(n416), .Z(n322) );
  NAND2_X1 U360 ( .A1(n48), .A2(n425), .ZN(n209) );
  INV_X1 U361 ( .A(n209), .ZN(n417) );
  MUX2_X1 U362 ( .A(\a[7][4] ), .B(data_in[4]), .S(n417), .Z(n326) );
  MUX2_X1 U363 ( .A(n34), .B(data_in[3]), .S(n417), .Z(n327) );
  MUX2_X1 U364 ( .A(\a[7][2] ), .B(data_in[2]), .S(n417), .Z(n328) );
  MUX2_X1 U365 ( .A(\a[7][1] ), .B(data_in[1]), .S(n417), .Z(n329) );
  MUX2_X1 U366 ( .A(\a[7][0] ), .B(data_in[0]), .S(n417), .Z(n330) );
  NAND2_X1 U367 ( .A1(n48), .A2(n78), .ZN(n32) );
  INV_X1 U368 ( .A(n32), .ZN(n418) );
  MUX2_X1 U369 ( .A(\a[6][4] ), .B(data_in[4]), .S(n418), .Z(n334) );
  MUX2_X1 U370 ( .A(\a[6][3] ), .B(data_in[3]), .S(n418), .Z(n335) );
  MUX2_X1 U371 ( .A(\a[6][2] ), .B(data_in[2]), .S(n418), .Z(n336) );
  MUX2_X1 U372 ( .A(n148), .B(data_in[1]), .S(n418), .Z(n337) );
  MUX2_X1 U373 ( .A(\a[6][0] ), .B(data_in[0]), .S(n418), .Z(n338) );
  NAND2_X1 U374 ( .A1(n48), .A2(n47), .ZN(n38) );
  INV_X1 U375 ( .A(n38), .ZN(n419) );
  MUX2_X1 U376 ( .A(\a[5][4] ), .B(data_in[4]), .S(n419), .Z(n342) );
  MUX2_X1 U377 ( .A(\a[5][3] ), .B(data_in[3]), .S(n419), .Z(n343) );
  MUX2_X1 U378 ( .A(\a[5][2] ), .B(data_in[2]), .S(n419), .Z(n344) );
  MUX2_X1 U379 ( .A(n96), .B(data_in[1]), .S(n419), .Z(n345) );
  MUX2_X1 U380 ( .A(\a[5][0] ), .B(data_in[0]), .S(n419), .Z(n346) );
  NAND2_X1 U381 ( .A1(n48), .A2(n58), .ZN(n49) );
  INV_X1 U382 ( .A(n49), .ZN(n420) );
  MUX2_X1 U383 ( .A(\a[4][4] ), .B(data_in[4]), .S(n420), .Z(n350) );
  MUX2_X1 U384 ( .A(n387), .B(data_in[3]), .S(n420), .Z(n351) );
  MUX2_X1 U385 ( .A(\a[4][2] ), .B(data_in[2]), .S(n420), .Z(n352) );
  MUX2_X1 U386 ( .A(n405), .B(data_in[1]), .S(n420), .Z(n353) );
  MUX2_X1 U387 ( .A(\a[4][0] ), .B(data_in[0]), .S(n420), .Z(n354) );
  NAND2_X1 U388 ( .A1(n68), .A2(n425), .ZN(n59) );
  INV_X1 U389 ( .A(n59), .ZN(n421) );
  MUX2_X1 U390 ( .A(\a[3][4] ), .B(data_in[4]), .S(n421), .Z(n358) );
  MUX2_X1 U391 ( .A(\a[3][3] ), .B(data_in[3]), .S(n421), .Z(n359) );
  MUX2_X1 U392 ( .A(\a[3][2] ), .B(data_in[2]), .S(n421), .Z(n360) );
  MUX2_X1 U393 ( .A(\a[3][1] ), .B(data_in[1]), .S(n421), .Z(n361) );
  MUX2_X1 U395 ( .A(\a[3][0] ), .B(data_in[0]), .S(n421), .Z(n362) );
  NAND2_X1 U396 ( .A1(n78), .A2(n68), .ZN(n69) );
  INV_X1 U397 ( .A(n69), .ZN(n422) );
  MUX2_X1 U398 ( .A(\a[2][4] ), .B(data_in[4]), .S(n422), .Z(n366) );
  MUX2_X1 U399 ( .A(\a[2][3] ), .B(data_in[3]), .S(n422), .Z(n367) );
  MUX2_X1 U400 ( .A(\a[2][2] ), .B(data_in[2]), .S(n422), .Z(n368) );
  MUX2_X1 U401 ( .A(n95), .B(data_in[1]), .S(n422), .Z(n369) );
  MUX2_X1 U402 ( .A(\a[2][0] ), .B(data_in[0]), .S(n422), .Z(n370) );
  NAND2_X1 U403 ( .A1(n47), .A2(n68), .ZN(n79) );
  INV_X1 U404 ( .A(n79), .ZN(n423) );
  MUX2_X1 U405 ( .A(\a[1][4] ), .B(data_in[4]), .S(n423), .Z(n374) );
  MUX2_X1 U406 ( .A(\a[1][3] ), .B(data_in[3]), .S(n423), .Z(n375) );
  MUX2_X1 U407 ( .A(\a[1][2] ), .B(data_in[2]), .S(n423), .Z(n376) );
  MUX2_X1 U408 ( .A(\a[1][1] ), .B(data_in[1]), .S(n423), .Z(n377) );
  MUX2_X1 U409 ( .A(\a[1][0] ), .B(data_in[0]), .S(n423), .Z(n378) );
  NAND2_X1 U410 ( .A1(n68), .A2(n58), .ZN(n88) );
  INV_X1 U411 ( .A(n88), .ZN(n424) );
  MUX2_X1 U412 ( .A(\a[0][4] ), .B(data_in[4]), .S(n424), .Z(n382) );
  MUX2_X1 U413 ( .A(\a[0][3] ), .B(data_in[3]), .S(n424), .Z(n383) );
  MUX2_X1 U414 ( .A(\a[0][2] ), .B(data_in[2]), .S(n424), .Z(n384) );
  MUX2_X1 U415 ( .A(\a[0][1] ), .B(data_in[1]), .S(n424), .Z(n385) );
  MUX2_X1 U416 ( .A(\a[0][0] ), .B(data_in[0]), .S(n424), .Z(n386) );
  INV_X1 U417 ( .A(data_in[3]), .ZN(n443) );
  INV_X1 U418 ( .A(data_in[4]), .ZN(n442) );
endmodule


module control_DELAY2 ( clk, reset, start, done, en_a, en_x, en_y, clr_addr_a, 
        clr_addr_x, clr_addr_y, clr_delay, of_a, of_x, of_y, of_delay );
  input clk, reset, start, of_a, of_x, of_y, of_delay;
  output done, en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay;
  wire   \in_state[1] , n1, n7, n8, n12, n14, n15, n16, n17, n18, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n2, n3, n4, n5,
         n6, n9, n10, n11, n13, n19, n20, n21, n22;
  wire   [1:0] out_state;

  DFF_X1 \in_state_reg[0]  ( .D(n63), .CK(clk), .QN(n8) );
  DFF_X1 \out_state_reg[0]  ( .D(n61), .CK(clk), .Q(out_state[0]), .QN(n14) );
  DFF_X1 \out_state_reg[1]  ( .D(n60), .CK(clk), .Q(out_state[1]), .QN(n12) );
  DFF_X1 done_reg ( .D(n59), .CK(clk), .Q(done), .QN(n1) );
  DFF_X1 en_a_reg ( .D(n58), .CK(clk), .Q(en_a) );
  DFF_X1 en_x_reg ( .D(n57), .CK(clk), .Q(en_x) );
  DFF_X1 clr_addr_a_reg ( .D(n55), .CK(clk), .Q(clr_addr_a), .QN(n16) );
  DFF_X1 clr_addr_x_reg ( .D(n54), .CK(clk), .Q(clr_addr_x), .QN(n17) );
  DFF_X1 clr_delay_reg ( .D(n6), .CK(clk), .Q(clr_delay) );
  NAND3_X1 U51 ( .A1(of_delay), .A2(n12), .A3(out_state[0]), .ZN(n35) );
  NAND3_X1 U52 ( .A1(n28), .A2(n21), .A3(n32), .ZN(n37) );
  NAND3_X1 U53 ( .A1(n12), .A2(n21), .A3(out_state[0]), .ZN(n33) );
  NAND3_X1 U54 ( .A1(n8), .A2(n14), .A3(n46), .ZN(n47) );
  NAND3_X1 U55 ( .A1(n49), .A2(n21), .A3(n32), .ZN(n50) );
  NAND3_X1 U56 ( .A1(n49), .A2(n21), .A3(n52), .ZN(n51) );
  DFF_X1 clr_addr_y_reg ( .D(n53), .CK(clk), .Q(clr_addr_y), .QN(n18) );
  DFF_X1 en_y_reg ( .D(n56), .CK(clk), .Q(en_y), .QN(n15) );
  DFF_X1 \in_state_reg[1]  ( .D(n62), .CK(clk), .Q(\in_state[1] ), .QN(n7) );
  INV_X1 U3 ( .A(n28), .ZN(n5) );
  INV_X1 U4 ( .A(n30), .ZN(n2) );
  OAI21_X1 U5 ( .B1(n22), .B2(n42), .A(n5), .ZN(n49) );
  OAI21_X1 U6 ( .B1(n40), .B2(n22), .A(n41), .ZN(n30) );
  AOI21_X1 U7 ( .B1(n4), .B2(of_x), .A(n3), .ZN(n40) );
  OAI21_X1 U8 ( .B1(n19), .B2(n43), .A(n41), .ZN(n28) );
  INV_X1 U9 ( .A(n43), .ZN(n4) );
  INV_X1 U10 ( .A(of_delay), .ZN(n20) );
  INV_X1 U11 ( .A(n42), .ZN(n3) );
  INV_X1 U12 ( .A(n26), .ZN(n11) );
  INV_X1 U13 ( .A(of_x), .ZN(n19) );
  OAI21_X1 U14 ( .B1(n34), .B2(n12), .A(n13), .ZN(n26) );
  INV_X1 U15 ( .A(n25), .ZN(n13) );
  NOR2_X1 U16 ( .A1(n8), .A2(\in_state[1] ), .ZN(n32) );
  AOI21_X1 U17 ( .B1(out_state[0]), .B2(out_state[1]), .A(reset), .ZN(n27) );
  AOI21_X1 U18 ( .B1(n32), .B2(of_a), .A(reset), .ZN(n41) );
  OAI22_X1 U19 ( .A1(n26), .A2(n15), .B1(n11), .B2(n33), .ZN(n56) );
  OAI22_X1 U20 ( .A1(n44), .A2(n1), .B1(n10), .B2(n33), .ZN(n59) );
  INV_X1 U21 ( .A(n44), .ZN(n10) );
  OAI21_X1 U22 ( .B1(n20), .B2(n14), .A(n27), .ZN(n44) );
  OAI22_X1 U23 ( .A1(n28), .A2(n17), .B1(n5), .B2(n29), .ZN(n54) );
  NOR2_X1 U24 ( .A1(n4), .A2(reset), .ZN(n29) );
  OAI22_X1 U25 ( .A1(n30), .A2(n16), .B1(n2), .B2(n31), .ZN(n55) );
  NOR2_X1 U26 ( .A1(n32), .A2(reset), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n26), .A2(n18), .B1(n11), .B2(n27), .ZN(n53) );
  NAND2_X1 U28 ( .A1(n8), .A2(n7), .ZN(n42) );
  NOR2_X1 U29 ( .A1(n19), .A2(n7), .ZN(n46) );
  NAND2_X1 U30 ( .A1(\in_state[1] ), .A2(n8), .ZN(n43) );
  AOI21_X1 U31 ( .B1(n9), .B2(n47), .A(reset), .ZN(n61) );
  INV_X1 U32 ( .A(n48), .ZN(n9) );
  AOI21_X1 U33 ( .B1(of_y), .B2(out_state[1]), .A(n14), .ZN(n48) );
  OAI21_X1 U34 ( .B1(n8), .B2(n49), .A(n51), .ZN(n63) );
  OAI21_X1 U35 ( .B1(n43), .B2(n22), .A(n42), .ZN(n52) );
  NAND2_X1 U36 ( .A1(n46), .A2(n8), .ZN(n24) );
  OAI21_X1 U37 ( .B1(n20), .B2(n33), .A(n45), .ZN(n60) );
  NAND4_X1 U38 ( .A1(out_state[1]), .A2(n34), .A3(n24), .A4(n21), .ZN(n45) );
  OAI21_X1 U39 ( .B1(n7), .B2(n49), .A(n50), .ZN(n62) );
  NAND2_X1 U40 ( .A1(n21), .A2(n35), .ZN(n25) );
  NAND2_X1 U41 ( .A1(of_y), .A2(out_state[0]), .ZN(n34) );
  NAND2_X1 U42 ( .A1(n36), .A2(n37), .ZN(n57) );
  NAND2_X1 U43 ( .A1(en_x), .A2(n5), .ZN(n36) );
  NAND2_X1 U44 ( .A1(n38), .A2(n39), .ZN(n58) );
  OAI211_X1 U45 ( .C1(n3), .C2(n4), .A(n30), .B(n21), .ZN(n39) );
  NAND2_X1 U46 ( .A1(en_a), .A2(n2), .ZN(n38) );
  INV_X1 U47 ( .A(n23), .ZN(n6) );
  AOI21_X1 U48 ( .B1(n24), .B2(clr_delay), .A(n25), .ZN(n23) );
  INV_X1 U49 ( .A(reset), .ZN(n21) );
  INV_X1 U50 ( .A(start), .ZN(n22) );
endmodule


module mvm4_part3 ( clk, reset, start, done, data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, start;
  output done;
  wire   en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay, of_a,
         of_x, of_y, of_delay;

  data_path_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_DELAY2 datapath ( 
        .clk(clk), .en_a(en_a), .en_x(en_x), .en_y(en_y), .clr_addr_a(
        clr_addr_a), .clr_addr_x(clr_addr_x), .clr_addr_y(clr_addr_y), 
        .clr_delay(clr_delay), .of_a(of_a), .of_x(of_x), .of_y(of_y), 
        .of_delay(of_delay), .data_in(data_in), .data_out(data_out) );
  control_DELAY2 ctrl ( .clk(clk), .reset(reset), .start(start), .done(done), 
        .en_a(en_a), .en_x(en_x), .en_y(en_y), .clr_addr_a(clr_addr_a), 
        .clr_addr_x(clr_addr_x), .clr_addr_y(clr_addr_y), .clr_delay(clr_delay), .of_a(of_a), .of_x(of_x), .of_y(of_y), .of_delay(of_delay) );
endmodule

