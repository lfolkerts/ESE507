
module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n67, n68, n69,
         n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86, n87, n90,
         n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n139,
         n140, n142, n143, n145, n146, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n227, n228, n229, n230, n232, n233, n234, n235, n236, n237, n238,
         n240, n241, n242, n243, n244, n245, n246, n247, n255, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n337, n338, n339, n340, n341, n342,
         n343;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n160), .B(n100), .CI(n153), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n330), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n111), .B(n162), .CI(n156), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n170), .B(n177), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n166), .B(n149), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  NOR2_X1 U249 ( .A1(n331), .A2(n55), .ZN(n50) );
  CLKBUF_X1 U250 ( .A(n246), .Z(n285) );
  CLKBUF_X1 U251 ( .A(n246), .Z(n286) );
  AOI21_X1 U252 ( .B1(n58), .B2(n50), .A(n51), .ZN(n287) );
  BUF_X2 U253 ( .A(n238), .Z(n337) );
  AND2_X1 U254 ( .A1(n102), .A2(n99), .ZN(n288) );
  OR2_X1 U255 ( .A1(n183), .A2(n151), .ZN(n289) );
  OAI21_X1 U256 ( .B1(n52), .B2(n56), .A(n53), .ZN(n290) );
  OAI21_X2 U257 ( .B1(n67), .B2(n69), .A(n68), .ZN(n302) );
  OR2_X1 U258 ( .A1(n125), .A2(n128), .ZN(n291) );
  CLKBUF_X1 U259 ( .A(n194), .Z(n292) );
  CLKBUF_X1 U260 ( .A(n343), .Z(n293) );
  BUF_X2 U261 ( .A(n227), .Z(n343) );
  CLKBUF_X1 U262 ( .A(n315), .Z(n294) );
  BUF_X2 U263 ( .A(n318), .Z(n295) );
  XNOR2_X1 U264 ( .A(n245), .B(a[6]), .ZN(n318) );
  AOI21_X1 U265 ( .B1(n333), .B2(n302), .A(n63), .ZN(n296) );
  XNOR2_X1 U266 ( .A(n245), .B(n321), .ZN(n229) );
  XOR2_X1 U267 ( .A(n246), .B(a[2]), .Z(n297) );
  BUF_X2 U268 ( .A(n247), .Z(n298) );
  CLKBUF_X1 U269 ( .A(n246), .Z(n299) );
  CLKBUF_X1 U270 ( .A(n247), .Z(n300) );
  XNOR2_X1 U271 ( .A(n115), .B(n301), .ZN(n113) );
  XNOR2_X1 U272 ( .A(n120), .B(n117), .ZN(n301) );
  CLKBUF_X1 U273 ( .A(n55), .Z(n303) );
  AOI21_X1 U274 ( .B1(n333), .B2(n302), .A(n63), .ZN(n304) );
  NAND2_X1 U275 ( .A1(n115), .A2(n120), .ZN(n305) );
  NAND2_X1 U276 ( .A1(n115), .A2(n117), .ZN(n306) );
  NAND2_X1 U277 ( .A1(n120), .A2(n117), .ZN(n307) );
  NAND3_X1 U278 ( .A1(n305), .A2(n306), .A3(n307), .ZN(n112) );
  BUF_X2 U279 ( .A(n244), .Z(n308) );
  XNOR2_X1 U280 ( .A(n247), .B(a[2]), .ZN(n309) );
  CLKBUF_X1 U281 ( .A(n314), .Z(n310) );
  CLKBUF_X1 U282 ( .A(n245), .Z(n311) );
  CLKBUF_X1 U283 ( .A(n56), .Z(n312) );
  CLKBUF_X1 U284 ( .A(n334), .Z(n313) );
  NAND2_X1 U285 ( .A1(n230), .A2(n309), .ZN(n314) );
  OAI21_X1 U286 ( .B1(n59), .B2(n61), .A(n60), .ZN(n315) );
  INV_X1 U287 ( .A(n288), .ZN(n316) );
  OR2_X2 U288 ( .A1(n317), .A2(n146), .ZN(n235) );
  XNOR2_X1 U289 ( .A(n247), .B(n146), .ZN(n317) );
  NAND2_X1 U290 ( .A1(n229), .A2(n237), .ZN(n319) );
  NAND2_X1 U291 ( .A1(n229), .A2(n237), .ZN(n233) );
  NAND2_X1 U292 ( .A1(n246), .A2(a[4]), .ZN(n322) );
  NAND2_X1 U293 ( .A1(n320), .A2(n321), .ZN(n323) );
  NAND2_X1 U294 ( .A1(n322), .A2(n323), .ZN(n237) );
  INV_X1 U295 ( .A(n246), .ZN(n320) );
  INV_X1 U296 ( .A(a[4]), .ZN(n321) );
  CLKBUF_X1 U297 ( .A(n246), .Z(n324) );
  CLKBUF_X1 U298 ( .A(n245), .Z(n325) );
  INV_X1 U299 ( .A(n45), .ZN(n326) );
  OAI21_X2 U300 ( .B1(n49), .B2(n37), .A(n38), .ZN(n36) );
  AOI21_X1 U301 ( .B1(n58), .B2(n50), .A(n51), .ZN(n327) );
  NOR2_X1 U302 ( .A1(n103), .A2(n106), .ZN(n328) );
  OAI21_X1 U303 ( .B1(n41), .B2(n47), .A(n42), .ZN(n329) );
  NAND2_X1 U304 ( .A1(n297), .A2(n309), .ZN(n234) );
  OAI22_X1 U305 ( .A1(n234), .A2(n203), .B1(n202), .B2(n337), .ZN(n330) );
  NOR2_X1 U306 ( .A1(n113), .A2(n118), .ZN(n331) );
  XNOR2_X1 U307 ( .A(n245), .B(a[6]), .ZN(n236) );
  INV_X1 U308 ( .A(n329), .ZN(n38) );
  INV_X1 U309 ( .A(n39), .ZN(n37) );
  XNOR2_X1 U310 ( .A(n48), .B(n5), .ZN(product[9]) );
  NAND2_X1 U311 ( .A1(n85), .A2(n326), .ZN(n5) );
  INV_X1 U312 ( .A(n46), .ZN(n85) );
  INV_X1 U313 ( .A(n47), .ZN(n45) );
  INV_X1 U314 ( .A(n77), .ZN(n75) );
  AOI21_X1 U315 ( .B1(n333), .B2(n302), .A(n63), .ZN(n61) );
  NOR2_X1 U316 ( .A1(n113), .A2(n118), .ZN(n52) );
  NOR2_X1 U317 ( .A1(n107), .A2(n112), .ZN(n46) );
  NAND2_X1 U318 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U319 ( .A(n71), .ZN(n91) );
  NAND2_X1 U320 ( .A1(n291), .A2(n60), .ZN(n8) );
  NAND2_X1 U321 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U322 ( .A(n20), .ZN(n81) );
  NAND2_X1 U323 ( .A1(n84), .A2(n42), .ZN(n4) );
  NAND2_X1 U324 ( .A1(n332), .A2(n30), .ZN(n2) );
  NAND2_X1 U325 ( .A1(n107), .A2(n112), .ZN(n47) );
  XOR2_X1 U326 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U327 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U328 ( .A(n67), .ZN(n90) );
  XNOR2_X1 U329 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U330 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U331 ( .B1(n57), .B2(n303), .A(n312), .ZN(n54) );
  XNOR2_X1 U332 ( .A(n9), .B(n302), .ZN(product[5]) );
  NAND2_X1 U333 ( .A1(n333), .A2(n65), .ZN(n9) );
  INV_X1 U334 ( .A(n70), .ZN(n69) );
  XNOR2_X1 U335 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U336 ( .A1(n335), .A2(n77), .ZN(n12) );
  XOR2_X1 U337 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U338 ( .A1(n87), .A2(n312), .ZN(n7) );
  INV_X1 U339 ( .A(n303), .ZN(n87) );
  INV_X1 U340 ( .A(n338), .ZN(n24) );
  OR2_X1 U341 ( .A1(n98), .A2(n97), .ZN(n332) );
  OR2_X1 U342 ( .A1(n129), .A2(n132), .ZN(n333) );
  NOR2_X1 U343 ( .A1(n119), .A2(n124), .ZN(n55) );
  INV_X1 U344 ( .A(n94), .ZN(n95) );
  NOR2_X1 U345 ( .A1(n125), .A2(n128), .ZN(n59) );
  NOR2_X1 U346 ( .A1(n96), .A2(n95), .ZN(n20) );
  NOR2_X1 U347 ( .A1(n133), .A2(n134), .ZN(n67) );
  NAND2_X1 U348 ( .A1(n119), .A2(n124), .ZN(n56) );
  OR2_X1 U349 ( .A1(n99), .A2(n102), .ZN(n334) );
  NAND2_X1 U350 ( .A1(n125), .A2(n128), .ZN(n60) );
  INV_X1 U351 ( .A(n80), .ZN(n78) );
  NAND2_X1 U352 ( .A1(n129), .A2(n132), .ZN(n65) );
  NAND2_X1 U353 ( .A1(n133), .A2(n134), .ZN(n68) );
  NAND2_X1 U354 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U355 ( .A1(n182), .A2(n175), .ZN(n335) );
  NAND2_X1 U356 ( .A1(n98), .A2(n97), .ZN(n30) );
  NAND2_X1 U357 ( .A1(n103), .A2(n106), .ZN(n42) );
  INV_X1 U358 ( .A(n14), .ZN(product[15]) );
  OR2_X1 U359 ( .A1(n343), .A2(n242), .ZN(n210) );
  AND2_X1 U360 ( .A1(n293), .A2(n140), .ZN(n167) );
  INV_X1 U361 ( .A(n100), .ZN(n101) );
  AND2_X1 U362 ( .A1(n343), .A2(n137), .ZN(n159) );
  INV_X1 U363 ( .A(n136), .ZN(n152) );
  OR2_X1 U364 ( .A1(n343), .A2(n240), .ZN(n192) );
  INV_X1 U365 ( .A(n139), .ZN(n160) );
  AND2_X1 U366 ( .A1(n289), .A2(n80), .ZN(product[1]) );
  OR2_X1 U367 ( .A1(n343), .A2(n241), .ZN(n201) );
  INV_X1 U368 ( .A(n146), .ZN(n255) );
  AND2_X1 U369 ( .A1(n293), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U370 ( .A(n247), .B(a[2]), .ZN(n238) );
  AOI21_X1 U371 ( .B1(n288), .B2(n332), .A(n28), .ZN(n338) );
  AOI21_X1 U372 ( .B1(n288), .B2(n332), .A(n28), .ZN(n26) );
  INV_X1 U373 ( .A(n30), .ZN(n28) );
  NAND2_X1 U374 ( .A1(n228), .A2(n318), .ZN(n339) );
  NAND2_X1 U375 ( .A1(n228), .A2(n295), .ZN(n340) );
  NAND2_X1 U376 ( .A1(n228), .A2(n236), .ZN(n232) );
  XOR2_X1 U377 ( .A(n244), .B(a[6]), .Z(n228) );
  INV_X1 U378 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U379 ( .A(n308), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U380 ( .A(n308), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U381 ( .A(n308), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U382 ( .A(n308), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U383 ( .A(n343), .B(n308), .ZN(n191) );
  NOR2_X1 U384 ( .A1(n46), .A2(n41), .ZN(n39) );
  INV_X1 U385 ( .A(n328), .ZN(n84) );
  NOR2_X1 U386 ( .A1(n103), .A2(n106), .ZN(n41) );
  INV_X1 U387 ( .A(n25), .ZN(n23) );
  NOR2_X1 U388 ( .A1(n25), .A2(n20), .ZN(n18) );
  NAND2_X1 U389 ( .A1(n113), .A2(n118), .ZN(n53) );
  XNOR2_X1 U390 ( .A(n308), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U391 ( .A(n246), .B(a[4]), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n246), .B(a[4]), .ZN(n342) );
  OAI22_X1 U393 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U394 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U395 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  OAI22_X1 U396 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U397 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U398 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OR2_X1 U399 ( .A1(n343), .A2(n243), .ZN(n219) );
  INV_X1 U400 ( .A(n145), .ZN(n176) );
  OR2_X1 U401 ( .A1(n169), .A2(n157), .ZN(n116) );
  XNOR2_X1 U402 ( .A(n169), .B(n157), .ZN(n117) );
  NAND2_X1 U403 ( .A1(n135), .A2(n150), .ZN(n72) );
  NOR2_X1 U404 ( .A1(n135), .A2(n150), .ZN(n71) );
  INV_X1 U405 ( .A(n110), .ZN(n111) );
  INV_X1 U406 ( .A(n142), .ZN(n168) );
  AND2_X1 U407 ( .A1(n343), .A2(n143), .ZN(n175) );
  XNOR2_X1 U408 ( .A(n308), .B(b[2]), .ZN(n189) );
  XOR2_X1 U409 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U410 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  AOI21_X1 U411 ( .B1(n335), .B2(n78), .A(n75), .ZN(n73) );
  NAND2_X1 U412 ( .A1(n183), .A2(n151), .ZN(n80) );
  INV_X1 U413 ( .A(n294), .ZN(n57) );
  OAI21_X1 U414 ( .B1(n59), .B2(n304), .A(n60), .ZN(n58) );
  OAI21_X1 U415 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  OAI21_X1 U416 ( .B1(n328), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U417 ( .A1(n334), .A2(n332), .ZN(n25) );
  NAND2_X1 U418 ( .A1(n313), .A2(n316), .ZN(n3) );
  XOR2_X1 U419 ( .A(n43), .B(n4), .Z(product[10]) );
  XOR2_X1 U420 ( .A(n8), .B(n296), .Z(product[6]) );
  OAI22_X1 U421 ( .A1(n319), .A2(n199), .B1(n198), .B2(n341), .ZN(n165) );
  OAI22_X1 U422 ( .A1(n319), .A2(n197), .B1(n196), .B2(n342), .ZN(n163) );
  OAI22_X1 U423 ( .A1(n319), .A2(n198), .B1(n197), .B2(n342), .ZN(n164) );
  INV_X1 U424 ( .A(n342), .ZN(n140) );
  OAI22_X1 U425 ( .A1(n319), .A2(n292), .B1(n193), .B2(n341), .ZN(n100) );
  OAI22_X1 U426 ( .A1(n193), .A2(n319), .B1(n193), .B2(n341), .ZN(n139) );
  XNOR2_X1 U427 ( .A(n299), .B(b[5]), .ZN(n204) );
  OAI22_X1 U428 ( .A1(n319), .A2(n196), .B1(n195), .B2(n342), .ZN(n162) );
  XNOR2_X1 U429 ( .A(n324), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U430 ( .A(n299), .B(b[4]), .ZN(n205) );
  OAI22_X1 U431 ( .A1(n233), .A2(n195), .B1(n194), .B2(n341), .ZN(n161) );
  OAI22_X1 U432 ( .A1(n233), .A2(n241), .B1(n201), .B2(n342), .ZN(n149) );
  OAI22_X1 U433 ( .A1(n233), .A2(n200), .B1(n199), .B2(n341), .ZN(n166) );
  XNOR2_X1 U434 ( .A(n324), .B(b[2]), .ZN(n207) );
  INV_X1 U435 ( .A(n324), .ZN(n242) );
  XNOR2_X1 U436 ( .A(n343), .B(n324), .ZN(n209) );
  XNOR2_X1 U437 ( .A(n286), .B(b[6]), .ZN(n203) );
  XOR2_X1 U438 ( .A(n246), .B(a[2]), .Z(n230) );
  XOR2_X1 U439 ( .A(n31), .B(n2), .Z(product[12]) );
  INV_X1 U440 ( .A(n331), .ZN(n86) );
  OAI22_X1 U441 ( .A1(n184), .A2(n339), .B1(n184), .B2(n295), .ZN(n136) );
  OAI21_X1 U442 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  OAI22_X1 U443 ( .A1(n340), .A2(n185), .B1(n184), .B2(n295), .ZN(n94) );
  OAI22_X1 U444 ( .A1(n339), .A2(n188), .B1(n187), .B2(n295), .ZN(n155) );
  OAI22_X1 U445 ( .A1(n340), .A2(n187), .B1(n186), .B2(n295), .ZN(n154) );
  OAI22_X1 U446 ( .A1(n340), .A2(n186), .B1(n185), .B2(n295), .ZN(n153) );
  OAI22_X1 U447 ( .A1(n339), .A2(n190), .B1(n189), .B2(n295), .ZN(n157) );
  INV_X1 U448 ( .A(n318), .ZN(n137) );
  OAI22_X1 U449 ( .A1(n339), .A2(n189), .B1(n188), .B2(n295), .ZN(n156) );
  OAI22_X1 U450 ( .A1(n232), .A2(n240), .B1(n192), .B2(n236), .ZN(n148) );
  OAI22_X1 U451 ( .A1(n232), .A2(n191), .B1(n190), .B2(n236), .ZN(n158) );
  XNOR2_X1 U452 ( .A(n325), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U453 ( .A(n311), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U454 ( .A(n325), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U455 ( .A(n325), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U456 ( .A(n311), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U457 ( .A(n325), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U458 ( .A(n343), .B(n311), .ZN(n200) );
  INV_X1 U459 ( .A(n245), .ZN(n241) );
  XOR2_X1 U460 ( .A(n22), .B(n1), .Z(product[13]) );
  INV_X1 U461 ( .A(n65), .ZN(n63) );
  OAI22_X1 U462 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  NAND2_X1 U463 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U464 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  AOI21_X1 U465 ( .B1(n50), .B2(n315), .A(n290), .ZN(n49) );
  OAI22_X1 U466 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  NAND2_X1 U467 ( .A1(n39), .A2(n18), .ZN(n16) );
  AOI21_X1 U468 ( .B1(n18), .B2(n40), .A(n19), .ZN(n17) );
  XNOR2_X1 U469 ( .A(n285), .B(b[7]), .ZN(n202) );
  AOI21_X1 U470 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  XNOR2_X1 U471 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U472 ( .A(n245), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U473 ( .A(n299), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U474 ( .A(n36), .B(n3), .ZN(product[11]) );
  AOI21_X1 U475 ( .B1(n36), .B2(n313), .A(n288), .ZN(n31) );
  AOI21_X1 U476 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U477 ( .B1(n327), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U478 ( .A(n287), .ZN(n48) );
  OAI22_X1 U479 ( .A1(n314), .A2(n204), .B1(n203), .B2(n337), .ZN(n169) );
  OAI22_X1 U480 ( .A1(n310), .A2(n207), .B1(n206), .B2(n337), .ZN(n172) );
  OAI22_X1 U481 ( .A1(n314), .A2(n206), .B1(n205), .B2(n337), .ZN(n171) );
  OAI22_X1 U482 ( .A1(n314), .A2(n205), .B1(n204), .B2(n337), .ZN(n170) );
  OAI22_X1 U483 ( .A1(n314), .A2(n208), .B1(n207), .B2(n337), .ZN(n173) );
  OAI22_X1 U484 ( .A1(n310), .A2(n242), .B1(n210), .B2(n337), .ZN(n150) );
  OAI22_X1 U485 ( .A1(n234), .A2(n203), .B1(n202), .B2(n337), .ZN(n110) );
  XNOR2_X1 U486 ( .A(n298), .B(b[5]), .ZN(n213) );
  OAI22_X1 U487 ( .A1(n202), .A2(n234), .B1(n202), .B2(n337), .ZN(n142) );
  XNOR2_X1 U488 ( .A(n298), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U489 ( .A(n300), .B(b[4]), .ZN(n214) );
  INV_X1 U490 ( .A(n337), .ZN(n143) );
  OAI22_X1 U491 ( .A1(n314), .A2(n209), .B1(n208), .B2(n337), .ZN(n174) );
  XNOR2_X1 U492 ( .A(n298), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U493 ( .A(n343), .B(n300), .ZN(n218) );
  XNOR2_X1 U494 ( .A(n298), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U495 ( .A(n300), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U496 ( .A(n300), .B(b[1]), .ZN(n217) );
  INV_X1 U497 ( .A(n298), .ZN(n243) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86,
         n87, n88, n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n142, n143, n145, n146, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n227, n228, n230, n231, n233, n234, n235, n236,
         n238, n240, n241, n242, n243, n244, n245, n246, n247, n255, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n322), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n111), .B(n162), .CI(n156), .CO(n108), .S(n109) );
  FA_X1 U117 ( .A(n120), .B(n117), .CI(n115), .CO(n112), .S(n113) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n170), .B(n177), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n171), .B(n159), .CI(n178), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  AND2_X1 U249 ( .A1(n102), .A2(n99), .ZN(n295) );
  BUF_X2 U250 ( .A(n246), .Z(n310) );
  INV_X1 U251 ( .A(n295), .ZN(n35) );
  OR2_X1 U252 ( .A1(n183), .A2(n151), .ZN(n285) );
  XNOR2_X1 U253 ( .A(n240), .B(n308), .ZN(n311) );
  CLKBUF_X1 U254 ( .A(n304), .Z(n286) );
  NOR2_X1 U255 ( .A1(n103), .A2(n106), .ZN(n287) );
  AOI21_X1 U256 ( .B1(n325), .B2(n66), .A(n63), .ZN(n288) );
  CLKBUF_X1 U257 ( .A(n330), .Z(n289) );
  BUF_X2 U258 ( .A(n238), .Z(n333) );
  OAI21_X1 U259 ( .B1(n288), .B2(n59), .A(n60), .ZN(n290) );
  INV_X1 U260 ( .A(n140), .ZN(n291) );
  CLKBUF_X1 U261 ( .A(n342), .Z(n292) );
  NOR2_X1 U262 ( .A1(n103), .A2(n106), .ZN(n41) );
  XNOR2_X1 U263 ( .A(n317), .B(b[7]), .ZN(n293) );
  CLKBUF_X1 U264 ( .A(n244), .Z(n294) );
  CLKBUF_X1 U265 ( .A(b[7]), .Z(n296) );
  OAI21_X1 U266 ( .B1(n41), .B2(n47), .A(n42), .ZN(n297) );
  CLKBUF_X1 U267 ( .A(n190), .Z(n298) );
  NAND2_X2 U268 ( .A1(n231), .A2(n255), .ZN(n299) );
  NAND2_X1 U269 ( .A1(n231), .A2(n255), .ZN(n235) );
  BUF_X2 U270 ( .A(n227), .Z(n342) );
  CLKBUF_X1 U271 ( .A(n55), .Z(n300) );
  CLKBUF_X1 U272 ( .A(n246), .Z(n301) );
  BUF_X2 U273 ( .A(n245), .Z(n312) );
  CLKBUF_X1 U274 ( .A(n246), .Z(n336) );
  XNOR2_X1 U275 ( .A(n245), .B(a[6]), .ZN(n302) );
  XNOR2_X1 U276 ( .A(n245), .B(a[6]), .ZN(n236) );
  BUF_X1 U277 ( .A(n319), .Z(n303) );
  NAND2_X1 U278 ( .A1(n326), .A2(n327), .ZN(n304) );
  NAND2_X1 U279 ( .A1(n326), .A2(n327), .ZN(n233) );
  NAND2_X1 U280 ( .A1(n228), .A2(n236), .ZN(n305) );
  NOR2_X1 U281 ( .A1(n323), .A2(n55), .ZN(n306) );
  CLKBUF_X1 U282 ( .A(n53), .Z(n307) );
  CLKBUF_X1 U283 ( .A(a[6]), .Z(n308) );
  CLKBUF_X2 U284 ( .A(n236), .Z(n324) );
  BUF_X2 U285 ( .A(n247), .Z(n317) );
  BUF_X2 U286 ( .A(n238), .Z(n332) );
  INV_X1 U287 ( .A(n240), .ZN(n309) );
  XNOR2_X2 U288 ( .A(n301), .B(a[4]), .ZN(n337) );
  NAND2_X1 U289 ( .A1(n247), .A2(n314), .ZN(n315) );
  NAND2_X1 U290 ( .A1(n313), .A2(n146), .ZN(n316) );
  NAND2_X1 U291 ( .A1(n315), .A2(n316), .ZN(n231) );
  INV_X1 U292 ( .A(n247), .ZN(n313) );
  INV_X1 U293 ( .A(n146), .ZN(n314) );
  CLKBUF_X1 U294 ( .A(n323), .Z(n318) );
  CLKBUF_X1 U295 ( .A(n245), .Z(n319) );
  AOI21_X1 U296 ( .B1(n306), .B2(n290), .A(n51), .ZN(n320) );
  AOI21_X1 U297 ( .B1(n50), .B2(n58), .A(n51), .ZN(n49) );
  AOI21_X1 U298 ( .B1(n295), .B2(n328), .A(n28), .ZN(n321) );
  OAI22_X1 U299 ( .A1(n340), .A2(n203), .B1(n202), .B2(n333), .ZN(n322) );
  NOR2_X1 U300 ( .A1(n118), .A2(n113), .ZN(n323) );
  NOR2_X1 U301 ( .A1(n119), .A2(n124), .ZN(n55) );
  NOR2_X1 U302 ( .A1(n125), .A2(n128), .ZN(n59) );
  OR2_X1 U303 ( .A1(n129), .A2(n132), .ZN(n325) );
  NAND2_X1 U304 ( .A1(n119), .A2(n124), .ZN(n56) );
  NOR2_X1 U305 ( .A1(n133), .A2(n134), .ZN(n67) );
  XOR2_X1 U306 ( .A(n245), .B(a[4]), .Z(n326) );
  XNOR2_X1 U307 ( .A(n246), .B(a[4]), .ZN(n327) );
  XNOR2_X1 U308 ( .A(n48), .B(n5), .ZN(product[9]) );
  NAND2_X1 U309 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U310 ( .A(n46), .ZN(n85) );
  INV_X1 U311 ( .A(n297), .ZN(n38) );
  INV_X1 U312 ( .A(n39), .ZN(n37) );
  INV_X1 U313 ( .A(n25), .ZN(n23) );
  INV_X1 U314 ( .A(n47), .ZN(n45) );
  NOR2_X1 U315 ( .A1(n113), .A2(n118), .ZN(n52) );
  NAND2_X1 U316 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U317 ( .A(n20), .ZN(n81) );
  NOR2_X1 U318 ( .A1(n107), .A2(n112), .ZN(n46) );
  NAND2_X1 U319 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U320 ( .A(n59), .ZN(n88) );
  NAND2_X1 U321 ( .A1(n84), .A2(n42), .ZN(n4) );
  NAND2_X1 U322 ( .A1(n328), .A2(n30), .ZN(n2) );
  NAND2_X1 U323 ( .A1(n107), .A2(n112), .ZN(n47) );
  AOI21_X1 U324 ( .B1(n295), .B2(n328), .A(n28), .ZN(n26) );
  INV_X1 U325 ( .A(n30), .ZN(n28) );
  NAND2_X1 U326 ( .A1(n325), .A2(n65), .ZN(n9) );
  XOR2_X1 U327 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U328 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U329 ( .A(n300), .ZN(n87) );
  XNOR2_X1 U330 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U331 ( .A1(n86), .A2(n307), .ZN(n6) );
  OAI21_X1 U332 ( .B1(n57), .B2(n300), .A(n56), .ZN(n54) );
  INV_X1 U333 ( .A(n318), .ZN(n86) );
  NOR2_X1 U334 ( .A1(n25), .A2(n20), .ZN(n18) );
  AOI21_X1 U335 ( .B1(n329), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U336 ( .A(n77), .ZN(n75) );
  XNOR2_X1 U337 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U338 ( .A1(n329), .A2(n77), .ZN(n12) );
  INV_X1 U339 ( .A(n65), .ZN(n63) );
  OR2_X1 U340 ( .A1(n98), .A2(n97), .ZN(n328) );
  OAI21_X1 U341 ( .B1(n61), .B2(n59), .A(n60), .ZN(n58) );
  NOR2_X1 U342 ( .A1(n96), .A2(n95), .ZN(n20) );
  INV_X1 U343 ( .A(n94), .ZN(n95) );
  INV_X1 U344 ( .A(n80), .ZN(n78) );
  OR2_X1 U345 ( .A1(n182), .A2(n175), .ZN(n329) );
  XOR2_X1 U346 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U347 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U348 ( .A(n67), .ZN(n90) );
  OR2_X1 U349 ( .A1(n99), .A2(n102), .ZN(n330) );
  OAI21_X1 U350 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  XOR2_X1 U351 ( .A(n11), .B(n73), .Z(product[3]) );
  NAND2_X1 U352 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U353 ( .A(n71), .ZN(n91) );
  NAND2_X1 U354 ( .A1(n125), .A2(n128), .ZN(n60) );
  NAND2_X1 U355 ( .A1(n96), .A2(n95), .ZN(n21) );
  NAND2_X1 U356 ( .A1(n103), .A2(n106), .ZN(n42) );
  INV_X1 U357 ( .A(n14), .ZN(product[15]) );
  OR2_X1 U358 ( .A1(n292), .A2(n242), .ZN(n210) );
  AND2_X1 U359 ( .A1(n342), .A2(n140), .ZN(n167) );
  OR2_X1 U360 ( .A1(n241), .A2(n342), .ZN(n201) );
  INV_X1 U361 ( .A(n100), .ZN(n101) );
  AND2_X1 U362 ( .A1(n342), .A2(n137), .ZN(n159) );
  INV_X1 U363 ( .A(n136), .ZN(n152) );
  NAND2_X1 U364 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U365 ( .A1(n342), .A2(n240), .ZN(n192) );
  AND2_X1 U366 ( .A1(n285), .A2(n80), .ZN(product[1]) );
  AND2_X1 U367 ( .A1(n292), .A2(n146), .ZN(product[0]) );
  NAND2_X1 U368 ( .A1(n98), .A2(n97), .ZN(n30) );
  XNOR2_X1 U369 ( .A(n247), .B(a[2]), .ZN(n238) );
  OAI22_X1 U370 ( .A1(n299), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U371 ( .A1(n299), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U372 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U373 ( .A1(n299), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OR2_X1 U374 ( .A1(n292), .A2(n243), .ZN(n219) );
  OR2_X1 U375 ( .A1(n169), .A2(n157), .ZN(n116) );
  XNOR2_X1 U376 ( .A(n169), .B(n157), .ZN(n117) );
  NAND2_X1 U377 ( .A1(n135), .A2(n150), .ZN(n72) );
  NOR2_X1 U378 ( .A1(n135), .A2(n150), .ZN(n71) );
  AND2_X1 U379 ( .A1(n342), .A2(n143), .ZN(n175) );
  INV_X1 U380 ( .A(n287), .ZN(n84) );
  OAI21_X1 U381 ( .B1(n287), .B2(n47), .A(n42), .ZN(n40) );
  NOR2_X1 U382 ( .A1(n46), .A2(n41), .ZN(n39) );
  INV_X1 U383 ( .A(n145), .ZN(n176) );
  NAND2_X1 U384 ( .A1(n182), .A2(n175), .ZN(n77) );
  NAND2_X1 U385 ( .A1(n311), .A2(n302), .ZN(n334) );
  NAND2_X1 U386 ( .A1(n324), .A2(n311), .ZN(n335) );
  XOR2_X1 U387 ( .A(n244), .B(a[6]), .Z(n228) );
  INV_X1 U388 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U389 ( .A(n309), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U390 ( .A(n309), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U391 ( .A(n309), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U392 ( .A(n294), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U393 ( .A(n342), .B(n294), .ZN(n191) );
  OAI22_X1 U394 ( .A1(n299), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OAI22_X1 U395 ( .A1(n293), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U396 ( .A1(n299), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U397 ( .A1(n299), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OAI22_X1 U398 ( .A1(n299), .A2(n212), .B1(n293), .B2(n255), .ZN(n177) );
  INV_X1 U399 ( .A(n142), .ZN(n168) );
  INV_X1 U400 ( .A(n319), .ZN(n241) );
  XNOR2_X1 U401 ( .A(n312), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U402 ( .A(n312), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U403 ( .A(n303), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U404 ( .A(n312), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U405 ( .A(n342), .B(n312), .ZN(n200) );
  NAND2_X1 U406 ( .A1(n289), .A2(n35), .ZN(n3) );
  NAND2_X1 U407 ( .A1(n330), .A2(n328), .ZN(n25) );
  INV_X1 U408 ( .A(n110), .ZN(n111) );
  OAI21_X1 U409 ( .B1(n67), .B2(n69), .A(n68), .ZN(n338) );
  OAI21_X1 U410 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  XNOR2_X1 U411 ( .A(n309), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U412 ( .A(n312), .B(b[6]), .ZN(n194) );
  INV_X1 U413 ( .A(n290), .ZN(n57) );
  OAI22_X1 U414 ( .A1(n184), .A2(n334), .B1(n184), .B2(n324), .ZN(n136) );
  OAI22_X1 U415 ( .A1(n335), .A2(n185), .B1(n184), .B2(n324), .ZN(n94) );
  OAI22_X1 U416 ( .A1(n334), .A2(n188), .B1(n187), .B2(n324), .ZN(n155) );
  OAI22_X1 U417 ( .A1(n335), .A2(n187), .B1(n186), .B2(n324), .ZN(n154) );
  OAI22_X1 U418 ( .A1(n335), .A2(n298), .B1(n189), .B2(n324), .ZN(n157) );
  OAI22_X1 U419 ( .A1(n334), .A2(n189), .B1(n188), .B2(n324), .ZN(n156) );
  INV_X1 U420 ( .A(n302), .ZN(n137) );
  OAI22_X1 U421 ( .A1(n305), .A2(n240), .B1(n192), .B2(n302), .ZN(n148) );
  OAI22_X1 U422 ( .A1(n305), .A2(n191), .B1(n190), .B2(n302), .ZN(n158) );
  AOI21_X1 U423 ( .B1(n325), .B2(n338), .A(n63), .ZN(n339) );
  NAND2_X1 U424 ( .A1(n238), .A2(n230), .ZN(n340) );
  AOI21_X1 U425 ( .B1(n325), .B2(n66), .A(n63), .ZN(n61) );
  NAND2_X1 U426 ( .A1(n230), .A2(n332), .ZN(n234) );
  INV_X1 U427 ( .A(n139), .ZN(n160) );
  OAI22_X1 U428 ( .A1(n334), .A2(n186), .B1(n185), .B2(n324), .ZN(n153) );
  INV_X1 U429 ( .A(n70), .ZN(n69) );
  XOR2_X1 U430 ( .A(n8), .B(n339), .Z(product[6]) );
  NAND2_X1 U431 ( .A1(n113), .A2(n118), .ZN(n53) );
  XNOR2_X1 U432 ( .A(n9), .B(n338), .ZN(product[5]) );
  NAND2_X1 U433 ( .A1(n129), .A2(n132), .ZN(n65) );
  XOR2_X1 U434 ( .A(n43), .B(n4), .Z(product[10]) );
  INV_X1 U435 ( .A(n321), .ZN(n24) );
  OAI21_X1 U436 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  XNOR2_X1 U437 ( .A(n309), .B(n296), .ZN(n184) );
  XNOR2_X1 U438 ( .A(n303), .B(n296), .ZN(n193) );
  OAI21_X1 U439 ( .B1(n320), .B2(n37), .A(n38), .ZN(n341) );
  XOR2_X1 U440 ( .A(n31), .B(n2), .Z(product[12]) );
  OAI21_X1 U441 ( .B1(n37), .B2(n49), .A(n38), .ZN(n36) );
  NAND2_X1 U442 ( .A1(n183), .A2(n151), .ZN(n80) );
  XNOR2_X1 U443 ( .A(n317), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U444 ( .A(n317), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U445 ( .A(n317), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U446 ( .A(n317), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U447 ( .A(n317), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U448 ( .A(n292), .B(n317), .ZN(n218) );
  XNOR2_X1 U449 ( .A(n317), .B(b[1]), .ZN(n217) );
  INV_X1 U450 ( .A(n317), .ZN(n243) );
  NAND2_X1 U451 ( .A1(n39), .A2(n18), .ZN(n16) );
  AOI21_X1 U452 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  OAI21_X1 U453 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  NOR2_X1 U454 ( .A1(n323), .A2(n55), .ZN(n50) );
  XOR2_X1 U455 ( .A(n22), .B(n1), .Z(product[13]) );
  OAI22_X1 U456 ( .A1(n286), .A2(n199), .B1(n198), .B2(n291), .ZN(n165) );
  OAI22_X1 U457 ( .A1(n304), .A2(n198), .B1(n197), .B2(n337), .ZN(n164) );
  OAI22_X1 U458 ( .A1(n304), .A2(n197), .B1(n196), .B2(n337), .ZN(n163) );
  OAI22_X1 U459 ( .A1(n304), .A2(n194), .B1(n193), .B2(n337), .ZN(n100) );
  OAI22_X1 U460 ( .A1(n304), .A2(n196), .B1(n195), .B2(n337), .ZN(n162) );
  INV_X1 U461 ( .A(n337), .ZN(n140) );
  OAI22_X1 U462 ( .A1(n193), .A2(n286), .B1(n193), .B2(n291), .ZN(n139) );
  OAI22_X1 U463 ( .A1(n233), .A2(n195), .B1(n194), .B2(n337), .ZN(n161) );
  XNOR2_X1 U464 ( .A(n310), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U465 ( .A(n310), .B(b[5]), .ZN(n204) );
  OAI22_X1 U466 ( .A1(n233), .A2(n241), .B1(n201), .B2(n337), .ZN(n149) );
  OAI22_X1 U467 ( .A1(n233), .A2(n200), .B1(n199), .B2(n327), .ZN(n166) );
  XNOR2_X1 U468 ( .A(n336), .B(b[2]), .ZN(n207) );
  INV_X1 U469 ( .A(n336), .ZN(n242) );
  XNOR2_X1 U470 ( .A(n310), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U471 ( .A(n292), .B(n310), .ZN(n209) );
  XNOR2_X1 U472 ( .A(n310), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U473 ( .A(n310), .B(b[7]), .ZN(n202) );
  XOR2_X1 U474 ( .A(n246), .B(a[2]), .Z(n230) );
  AOI21_X1 U475 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  XNOR2_X1 U476 ( .A(n336), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U477 ( .A(n309), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U478 ( .A(n312), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U479 ( .A(n317), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U480 ( .A(n341), .B(n3), .ZN(product[11]) );
  AOI21_X1 U481 ( .B1(n36), .B2(n289), .A(n295), .ZN(n31) );
  AOI21_X1 U482 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U483 ( .B1(n49), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U484 ( .A(n320), .ZN(n48) );
  OAI22_X1 U485 ( .A1(n234), .A2(n204), .B1(n203), .B2(n333), .ZN(n169) );
  OAI22_X1 U486 ( .A1(n234), .A2(n207), .B1(n206), .B2(n332), .ZN(n172) );
  OAI22_X1 U487 ( .A1(n340), .A2(n206), .B1(n205), .B2(n332), .ZN(n171) );
  OAI22_X1 U488 ( .A1(n340), .A2(n205), .B1(n204), .B2(n333), .ZN(n170) );
  OAI22_X1 U489 ( .A1(n234), .A2(n208), .B1(n207), .B2(n333), .ZN(n173) );
  OAI22_X1 U490 ( .A1(n234), .A2(n242), .B1(n210), .B2(n333), .ZN(n150) );
  OAI22_X1 U491 ( .A1(n340), .A2(n203), .B1(n202), .B2(n333), .ZN(n110) );
  OAI22_X1 U492 ( .A1(n340), .A2(n202), .B1(n202), .B2(n332), .ZN(n142) );
  INV_X1 U493 ( .A(n333), .ZN(n143) );
  OAI22_X1 U494 ( .A1(n234), .A2(n209), .B1(n208), .B2(n332), .ZN(n174) );
  INV_X2 U495 ( .A(n146), .ZN(n255) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n33, n35, n36, n37,
         n38, n39, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n75, n77, n78, n80, n81, n85, n86, n87, n88, n90,
         n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n139, n140,
         n142, n143, n145, n146, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n240, n241, n242, n243, n244, n245, n246, n247, n255, n285, n286,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n331), .B(n161), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n156), .B(n162), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n177), .B(n170), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n171), .B(n159), .CI(n178), .CO(n126), .S(n127) );
  HA_X1 U127 ( .A(n166), .B(n149), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n181), .B(n174), .CO(n134), .S(n135) );
  XNOR2_X1 U249 ( .A(n169), .B(n157), .ZN(n117) );
  NAND3_X1 U250 ( .A1(n324), .A2(n325), .A3(n326), .ZN(n112) );
  OR2_X1 U251 ( .A1(n99), .A2(n102), .ZN(n334) );
  OR2_X1 U252 ( .A1(n98), .A2(n97), .ZN(n285) );
  OR2_X1 U253 ( .A1(n129), .A2(n132), .ZN(n286) );
  AND3_X1 U254 ( .A1(n308), .A2(n307), .A3(n309), .ZN(product[15]) );
  AND2_X1 U255 ( .A1(n335), .A2(n80), .ZN(product[1]) );
  CLKBUF_X1 U256 ( .A(n36), .Z(n289) );
  OAI21_X1 U257 ( .B1(n49), .B2(n37), .A(n38), .ZN(n36) );
  CLKBUF_X1 U258 ( .A(n131), .Z(n290) );
  CLKBUF_X1 U259 ( .A(n246), .Z(n291) );
  CLKBUF_X1 U260 ( .A(n320), .Z(n292) );
  OAI21_X1 U261 ( .B1(n329), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U262 ( .A(n146), .ZN(n293) );
  BUF_X1 U263 ( .A(n323), .Z(n294) );
  BUF_X2 U264 ( .A(n238), .Z(n340) );
  XNOR2_X1 U265 ( .A(n321), .B(a[2]), .ZN(n295) );
  XOR2_X1 U266 ( .A(n338), .B(a[4]), .Z(n296) );
  CLKBUF_X3 U267 ( .A(n245), .Z(n338) );
  NOR2_X1 U268 ( .A1(n25), .A2(n20), .ZN(n297) );
  INV_X2 U269 ( .A(n240), .ZN(n298) );
  BUF_X2 U270 ( .A(n338), .Z(n337) );
  XNOR2_X1 U271 ( .A(n22), .B(n299), .ZN(product[13]) );
  AND2_X1 U272 ( .A1(n81), .A2(n21), .ZN(n299) );
  CLKBUF_X1 U273 ( .A(n246), .Z(n300) );
  XNOR2_X1 U274 ( .A(n336), .B(a[6]), .ZN(n301) );
  CLKBUF_X1 U275 ( .A(n245), .Z(n336) );
  OR2_X1 U276 ( .A1(n103), .A2(n106), .ZN(n302) );
  XNOR2_X1 U277 ( .A(n115), .B(n315), .ZN(n303) );
  XNOR2_X1 U278 ( .A(n31), .B(n304), .ZN(product[12]) );
  AND2_X1 U279 ( .A1(n285), .A2(n30), .ZN(n304) );
  OAI21_X2 U280 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  NOR2_X1 U281 ( .A1(n103), .A2(n106), .ZN(n41) );
  OAI21_X1 U282 ( .B1(n52), .B2(n56), .A(n53), .ZN(n305) );
  XOR2_X1 U283 ( .A(n152), .B(n94), .Z(n306) );
  XOR2_X1 U284 ( .A(n15), .B(n306), .Z(product[14]) );
  NAND2_X1 U285 ( .A1(n15), .A2(n152), .ZN(n307) );
  NAND2_X1 U286 ( .A1(n15), .A2(n94), .ZN(n308) );
  NAND2_X1 U287 ( .A1(n152), .A2(n94), .ZN(n309) );
  BUF_X1 U288 ( .A(n247), .Z(n323) );
  OAI21_X1 U289 ( .B1(n41), .B2(n47), .A(n42), .ZN(n310) );
  NOR2_X1 U290 ( .A1(n125), .A2(n128), .ZN(n311) );
  INV_X1 U291 ( .A(n236), .ZN(n312) );
  INV_X1 U292 ( .A(n312), .ZN(n313) );
  NOR2_X1 U293 ( .A1(n125), .A2(n128), .ZN(n59) );
  XNOR2_X1 U294 ( .A(n323), .B(n293), .ZN(n231) );
  XNOR2_X1 U295 ( .A(n131), .B(n314), .ZN(n129) );
  XNOR2_X1 U296 ( .A(n172), .B(n179), .ZN(n314) );
  XNOR2_X1 U297 ( .A(n115), .B(n315), .ZN(n113) );
  XNOR2_X1 U298 ( .A(n120), .B(n117), .ZN(n315) );
  AOI21_X1 U299 ( .B1(n286), .B2(n66), .A(n63), .ZN(n316) );
  BUF_X1 U300 ( .A(n247), .Z(n321) );
  AOI21_X1 U301 ( .B1(n286), .B2(n66), .A(n63), .ZN(n61) );
  NAND2_X1 U302 ( .A1(n290), .A2(n172), .ZN(n317) );
  NAND2_X1 U303 ( .A1(n290), .A2(n179), .ZN(n318) );
  NAND2_X1 U304 ( .A1(n172), .A2(n179), .ZN(n319) );
  NAND3_X1 U305 ( .A1(n317), .A2(n318), .A3(n319), .ZN(n128) );
  NAND2_X1 U306 ( .A1(n230), .A2(n295), .ZN(n320) );
  CLKBUF_X1 U307 ( .A(n247), .Z(n322) );
  NAND2_X1 U308 ( .A1(n295), .A2(n230), .ZN(n234) );
  NAND2_X1 U309 ( .A1(n115), .A2(n120), .ZN(n324) );
  NAND2_X1 U310 ( .A1(n115), .A2(n117), .ZN(n325) );
  NAND2_X1 U311 ( .A1(n120), .A2(n117), .ZN(n326) );
  CLKBUF_X1 U312 ( .A(n238), .Z(n339) );
  XNOR2_X1 U313 ( .A(n246), .B(a[4]), .ZN(n327) );
  OAI21_X1 U314 ( .B1(n311), .B2(n61), .A(n60), .ZN(n328) );
  AOI21_X1 U315 ( .B1(n58), .B2(n50), .A(n305), .ZN(n329) );
  AOI21_X1 U316 ( .B1(n33), .B2(n285), .A(n28), .ZN(n330) );
  OAI22_X1 U317 ( .A1(n234), .A2(n203), .B1(n202), .B2(n340), .ZN(n331) );
  NOR2_X1 U318 ( .A1(n303), .A2(n118), .ZN(n332) );
  NOR2_X1 U319 ( .A1(n119), .A2(n124), .ZN(n55) );
  NAND2_X1 U320 ( .A1(n119), .A2(n124), .ZN(n56) );
  INV_X1 U321 ( .A(n310), .ZN(n38) );
  INV_X1 U322 ( .A(n39), .ZN(n37) );
  NAND2_X1 U323 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U324 ( .A(n328), .ZN(n57) );
  INV_X1 U325 ( .A(n46), .ZN(n85) );
  INV_X1 U326 ( .A(n47), .ZN(n45) );
  INV_X1 U327 ( .A(n25), .ZN(n23) );
  INV_X1 U328 ( .A(n30), .ZN(n28) );
  NOR2_X1 U329 ( .A1(n107), .A2(n112), .ZN(n46) );
  INV_X1 U330 ( .A(n65), .ZN(n63) );
  AOI21_X1 U331 ( .B1(n333), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U332 ( .A(n77), .ZN(n75) );
  NOR2_X1 U333 ( .A1(n113), .A2(n118), .ZN(n52) );
  NAND2_X1 U334 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U335 ( .A(n311), .ZN(n88) );
  INV_X1 U336 ( .A(n20), .ZN(n81) );
  NAND2_X1 U337 ( .A1(n286), .A2(n65), .ZN(n9) );
  XOR2_X1 U338 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U339 ( .A1(n302), .A2(n42), .ZN(n4) );
  XNOR2_X1 U340 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U341 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U342 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  XNOR2_X1 U343 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U344 ( .A1(n333), .A2(n77), .ZN(n12) );
  NOR2_X1 U345 ( .A1(n46), .A2(n41), .ZN(n39) );
  XOR2_X1 U346 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U347 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U348 ( .A(n55), .ZN(n87) );
  NAND2_X1 U349 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U350 ( .A(n71), .ZN(n91) );
  OR2_X1 U351 ( .A1(n169), .A2(n157), .ZN(n116) );
  INV_X1 U352 ( .A(n94), .ZN(n95) );
  NOR2_X1 U353 ( .A1(n96), .A2(n95), .ZN(n20) );
  XOR2_X1 U354 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U355 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U356 ( .A(n67), .ZN(n90) );
  OR2_X1 U357 ( .A1(n182), .A2(n175), .ZN(n333) );
  INV_X1 U358 ( .A(n70), .ZN(n69) );
  NAND2_X1 U359 ( .A1(n96), .A2(n95), .ZN(n21) );
  NAND2_X1 U360 ( .A1(n103), .A2(n106), .ZN(n42) );
  NAND2_X1 U361 ( .A1(n125), .A2(n128), .ZN(n60) );
  AND2_X1 U362 ( .A1(n227), .A2(n143), .ZN(n175) );
  OR2_X1 U363 ( .A1(n183), .A2(n151), .ZN(n335) );
  OR2_X1 U364 ( .A1(n227), .A2(n243), .ZN(n219) );
  OAI22_X1 U365 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  AND2_X1 U366 ( .A1(n227), .A2(n140), .ZN(n167) );
  OAI22_X1 U367 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OR2_X1 U368 ( .A1(n227), .A2(n241), .ZN(n201) );
  OAI22_X1 U369 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  NOR2_X1 U370 ( .A1(n133), .A2(n134), .ZN(n67) );
  INV_X1 U371 ( .A(n139), .ZN(n160) );
  OAI22_X1 U372 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  AND2_X1 U373 ( .A1(n227), .A2(n312), .ZN(n159) );
  INV_X1 U374 ( .A(n100), .ZN(n101) );
  INV_X1 U375 ( .A(n136), .ZN(n152) );
  NAND2_X1 U376 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U377 ( .A1(n227), .A2(n240), .ZN(n192) );
  OR2_X1 U378 ( .A1(n227), .A2(n242), .ZN(n210) );
  OAI22_X1 U379 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  AND2_X1 U380 ( .A1(n227), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U381 ( .A(n246), .B(a[4]), .ZN(n237) );
  XNOR2_X1 U382 ( .A(n321), .B(a[2]), .ZN(n238) );
  NAND2_X1 U383 ( .A1(n303), .A2(n118), .ZN(n53) );
  AOI21_X1 U384 ( .B1(n33), .B2(n285), .A(n28), .ZN(n26) );
  NAND2_X1 U385 ( .A1(n334), .A2(n285), .ZN(n25) );
  OAI21_X1 U386 ( .B1(n59), .B2(n316), .A(n60), .ZN(n58) );
  NAND2_X1 U387 ( .A1(n107), .A2(n112), .ZN(n47) );
  INV_X1 U388 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U389 ( .A(n227), .B(n244), .ZN(n191) );
  XNOR2_X1 U390 ( .A(n298), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U391 ( .A(n298), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U392 ( .A(n298), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U393 ( .A(n298), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U394 ( .A(n298), .B(b[7]), .ZN(n184) );
  INV_X1 U395 ( .A(n142), .ZN(n168) );
  XOR2_X1 U396 ( .A(n244), .B(a[6]), .Z(n228) );
  INV_X1 U397 ( .A(n110), .ZN(n111) );
  INV_X1 U398 ( .A(n35), .ZN(n33) );
  NAND2_X1 U399 ( .A1(n334), .A2(n35), .ZN(n3) );
  XNOR2_X1 U400 ( .A(n9), .B(n66), .ZN(product[5]) );
  NAND2_X1 U401 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U402 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  INV_X1 U403 ( .A(n145), .ZN(n176) );
  XNOR2_X1 U404 ( .A(n336), .B(a[6]), .ZN(n236) );
  XOR2_X1 U405 ( .A(n11), .B(n73), .Z(product[3]) );
  INV_X1 U406 ( .A(n80), .ZN(n78) );
  NAND2_X1 U407 ( .A1(n296), .A2(n237), .ZN(n341) );
  NAND2_X1 U408 ( .A1(n296), .A2(n327), .ZN(n342) );
  NAND2_X1 U409 ( .A1(n229), .A2(n237), .ZN(n233) );
  NOR2_X1 U410 ( .A1(n25), .A2(n20), .ZN(n18) );
  OAI22_X1 U411 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U412 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  NAND2_X1 U413 ( .A1(n129), .A2(n132), .ZN(n65) );
  NOR2_X1 U414 ( .A1(n135), .A2(n150), .ZN(n71) );
  INV_X1 U415 ( .A(n330), .ZN(n24) );
  OAI21_X1 U416 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U417 ( .A1(n98), .A2(n97), .ZN(n30) );
  XNOR2_X1 U418 ( .A(n298), .B(b[2]), .ZN(n189) );
  NAND2_X2 U419 ( .A1(n231), .A2(n255), .ZN(n235) );
  NAND2_X1 U420 ( .A1(n183), .A2(n151), .ZN(n80) );
  OAI21_X1 U421 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  OAI22_X1 U422 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  AOI21_X1 U423 ( .B1(n50), .B2(n328), .A(n51), .ZN(n49) );
  INV_X1 U424 ( .A(n332), .ZN(n86) );
  NOR2_X1 U425 ( .A1(n332), .A2(n55), .ZN(n50) );
  OAI22_X1 U426 ( .A1(n184), .A2(n232), .B1(n184), .B2(n313), .ZN(n136) );
  OAI21_X1 U427 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  OAI22_X1 U428 ( .A1(n232), .A2(n185), .B1(n184), .B2(n313), .ZN(n94) );
  OAI22_X1 U429 ( .A1(n232), .A2(n188), .B1(n187), .B2(n313), .ZN(n155) );
  OAI22_X1 U430 ( .A1(n232), .A2(n187), .B1(n186), .B2(n313), .ZN(n154) );
  OAI22_X1 U431 ( .A1(n232), .A2(n186), .B1(n185), .B2(n313), .ZN(n153) );
  OAI22_X1 U432 ( .A1(n232), .A2(n190), .B1(n189), .B2(n236), .ZN(n157) );
  OAI22_X1 U433 ( .A1(n232), .A2(n189), .B1(n236), .B2(n188), .ZN(n156) );
  OAI22_X1 U434 ( .A1(n232), .A2(n240), .B1(n192), .B2(n236), .ZN(n148) );
  OAI22_X1 U435 ( .A1(n232), .A2(n191), .B1(n190), .B2(n236), .ZN(n158) );
  XNOR2_X1 U436 ( .A(n337), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U437 ( .A(n337), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U438 ( .A(n338), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U439 ( .A(n337), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U440 ( .A(n227), .B(n337), .ZN(n200) );
  XNOR2_X1 U441 ( .A(n338), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U442 ( .A(b[7]), .B(n338), .ZN(n193) );
  INV_X1 U443 ( .A(n337), .ZN(n241) );
  NAND2_X2 U444 ( .A1(n228), .A2(n301), .ZN(n232) );
  XOR2_X1 U445 ( .A(n338), .B(a[4]), .Z(n229) );
  NAND2_X1 U446 ( .A1(n39), .A2(n297), .ZN(n16) );
  AOI21_X1 U447 ( .B1(n310), .B2(n18), .A(n19), .ZN(n17) );
  NAND2_X1 U448 ( .A1(n99), .A2(n102), .ZN(n35) );
  NAND2_X1 U449 ( .A1(n135), .A2(n150), .ZN(n72) );
  XNOR2_X1 U450 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U451 ( .A(n8), .B(n316), .Z(product[6]) );
  AOI21_X1 U452 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  OAI22_X1 U453 ( .A1(n341), .A2(n199), .B1(n198), .B2(n237), .ZN(n165) );
  OAI22_X1 U454 ( .A1(n342), .A2(n197), .B1(n196), .B2(n327), .ZN(n163) );
  OAI22_X1 U455 ( .A1(n342), .A2(n194), .B1(n193), .B2(n237), .ZN(n100) );
  OAI22_X1 U456 ( .A1(n342), .A2(n196), .B1(n195), .B2(n237), .ZN(n162) );
  OAI22_X1 U457 ( .A1(n233), .A2(n198), .B1(n197), .B2(n327), .ZN(n164) );
  OAI22_X1 U458 ( .A1(n193), .A2(n341), .B1(n193), .B2(n327), .ZN(n139) );
  OAI22_X1 U459 ( .A1(n195), .A2(n233), .B1(n194), .B2(n237), .ZN(n161) );
  INV_X1 U460 ( .A(n327), .ZN(n140) );
  OAI22_X1 U461 ( .A1(n233), .A2(n241), .B1(n201), .B2(n327), .ZN(n149) );
  XNOR2_X1 U462 ( .A(n300), .B(b[3]), .ZN(n206) );
  OAI22_X1 U463 ( .A1(n341), .A2(n200), .B1(n199), .B2(n327), .ZN(n166) );
  XNOR2_X1 U464 ( .A(n291), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U465 ( .A(n300), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U466 ( .A(n291), .B(b[5]), .ZN(n204) );
  INV_X1 U467 ( .A(n300), .ZN(n242) );
  XNOR2_X1 U468 ( .A(n291), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U469 ( .A(n246), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U470 ( .A(n227), .B(n300), .ZN(n209) );
  XOR2_X1 U471 ( .A(n246), .B(a[2]), .Z(n230) );
  XNOR2_X1 U472 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U473 ( .A(n338), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U474 ( .A(n300), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U475 ( .A(n289), .B(n3), .ZN(product[11]) );
  AOI21_X1 U476 ( .B1(n36), .B2(n334), .A(n33), .ZN(n31) );
  AOI21_X1 U477 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U478 ( .A(n329), .ZN(n48) );
  OAI22_X1 U479 ( .A1(n320), .A2(n204), .B1(n203), .B2(n339), .ZN(n169) );
  OAI22_X1 U480 ( .A1(n292), .A2(n207), .B1(n206), .B2(n339), .ZN(n172) );
  OAI22_X1 U481 ( .A1(n320), .A2(n206), .B1(n205), .B2(n340), .ZN(n171) );
  OAI22_X1 U482 ( .A1(n320), .A2(n205), .B1(n204), .B2(n340), .ZN(n170) );
  OAI22_X1 U483 ( .A1(n320), .A2(n208), .B1(n207), .B2(n339), .ZN(n173) );
  OAI22_X1 U484 ( .A1(n292), .A2(n242), .B1(n210), .B2(n339), .ZN(n150) );
  OAI22_X1 U485 ( .A1(n234), .A2(n203), .B1(n202), .B2(n340), .ZN(n110) );
  XNOR2_X1 U486 ( .A(n294), .B(b[5]), .ZN(n213) );
  OAI22_X1 U487 ( .A1(n202), .A2(n234), .B1(n202), .B2(n340), .ZN(n142) );
  XNOR2_X1 U488 ( .A(n294), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U489 ( .A(n322), .B(b[4]), .ZN(n214) );
  INV_X1 U490 ( .A(n340), .ZN(n143) );
  OAI22_X1 U491 ( .A1(n234), .A2(n209), .B1(n208), .B2(n339), .ZN(n174) );
  XNOR2_X1 U492 ( .A(n294), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U493 ( .A(n227), .B(n322), .ZN(n218) );
  XNOR2_X1 U494 ( .A(n322), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U495 ( .A(n322), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U496 ( .A(n322), .B(b[1]), .ZN(n217) );
  INV_X1 U497 ( .A(n323), .ZN(n243) );
  INV_X2 U498 ( .A(n146), .ZN(n255) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n24, n25, n26, n28, n30, n31, n36, n37, n38, n39,
         n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86, n87, n88, n90,
         n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n139, n140,
         n142, n143, n145, n146, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n227,
         n228, n230, n231, n232, n233, n234, n235, n236, n237, n238, n240,
         n241, n242, n243, n244, n245, n246, n247, n255, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n287), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n156), .B(n162), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n177), .B(n164), .CI(n170), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n166), .B(n149), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  CLKBUF_X3 U249 ( .A(n245), .Z(n325) );
  XNOR2_X1 U250 ( .A(n169), .B(n157), .ZN(n117) );
  AND2_X1 U251 ( .A1(n102), .A2(n99), .ZN(n285) );
  OR2_X1 U252 ( .A1(n183), .A2(n289), .ZN(n286) );
  OAI22_X1 U253 ( .A1(n234), .A2(n203), .B1(n202), .B2(n320), .ZN(n287) );
  OAI21_X1 U254 ( .B1(n52), .B2(n56), .A(n53), .ZN(n288) );
  OR2_X1 U255 ( .A1(n102), .A2(n99), .ZN(n335) );
  CLKBUF_X1 U256 ( .A(n151), .Z(n289) );
  OAI22_X1 U257 ( .A1(n328), .A2(n194), .B1(n193), .B2(n340), .ZN(n290) );
  CLKBUF_X1 U258 ( .A(n247), .Z(n316) );
  BUF_X1 U259 ( .A(n320), .Z(n291) );
  CLKBUF_X1 U260 ( .A(n328), .Z(n292) );
  CLKBUF_X1 U261 ( .A(n246), .Z(n293) );
  OAI21_X1 U262 ( .B1(n302), .B2(n47), .A(n42), .ZN(n294) );
  AOI21_X1 U263 ( .B1(n338), .B2(n66), .A(n63), .ZN(n295) );
  AND2_X1 U264 ( .A1(n335), .A2(n336), .ZN(n296) );
  XOR2_X1 U265 ( .A(n101), .B(n154), .Z(n297) );
  XOR2_X1 U266 ( .A(n104), .B(n297), .Z(n99) );
  NAND2_X1 U267 ( .A1(n104), .A2(n101), .ZN(n298) );
  NAND2_X1 U268 ( .A1(n104), .A2(n154), .ZN(n299) );
  NAND2_X1 U269 ( .A1(n101), .A2(n154), .ZN(n300) );
  NAND3_X1 U270 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n98) );
  OR2_X2 U271 ( .A1(n98), .A2(n97), .ZN(n336) );
  INV_X1 U272 ( .A(n303), .ZN(n301) );
  NOR2_X1 U273 ( .A1(n103), .A2(n106), .ZN(n302) );
  CLKBUF_X1 U274 ( .A(n285), .Z(n303) );
  BUF_X2 U275 ( .A(n305), .Z(n304) );
  XNOR2_X1 U276 ( .A(n246), .B(a[4]), .ZN(n305) );
  BUF_X1 U277 ( .A(n237), .Z(n340) );
  AOI21_X1 U278 ( .B1(n50), .B2(n307), .A(n288), .ZN(n306) );
  OAI21_X1 U279 ( .B1(n59), .B2(n295), .A(n60), .ZN(n307) );
  AOI21_X1 U280 ( .B1(n50), .B2(n58), .A(n51), .ZN(n49) );
  XNOR2_X1 U281 ( .A(n22), .B(n308), .ZN(product[13]) );
  AND2_X1 U282 ( .A1(n81), .A2(n21), .ZN(n308) );
  XNOR2_X1 U283 ( .A(n31), .B(n309), .ZN(product[12]) );
  AND2_X1 U284 ( .A1(n336), .A2(n30), .ZN(n309) );
  XNOR2_X1 U285 ( .A(n115), .B(n310), .ZN(n113) );
  XNOR2_X1 U286 ( .A(n120), .B(n117), .ZN(n310) );
  OAI21_X1 U287 ( .B1(n67), .B2(n69), .A(n68), .ZN(n311) );
  NAND2_X1 U288 ( .A1(n246), .A2(n313), .ZN(n314) );
  NAND2_X1 U289 ( .A1(n312), .A2(a[2]), .ZN(n315) );
  NAND2_X1 U290 ( .A1(n314), .A2(n315), .ZN(n230) );
  INV_X1 U291 ( .A(n246), .ZN(n312) );
  INV_X1 U292 ( .A(a[2]), .ZN(n313) );
  CLKBUF_X1 U293 ( .A(n295), .Z(n317) );
  CLKBUF_X1 U294 ( .A(n246), .Z(n318) );
  NAND2_X1 U295 ( .A1(n230), .A2(n320), .ZN(n319) );
  XNOR2_X1 U296 ( .A(n247), .B(a[2]), .ZN(n320) );
  CLKBUF_X1 U297 ( .A(n59), .Z(n321) );
  NAND2_X1 U298 ( .A1(n115), .A2(n120), .ZN(n322) );
  NAND2_X1 U299 ( .A1(n115), .A2(n117), .ZN(n323) );
  NAND2_X1 U300 ( .A1(n120), .A2(n117), .ZN(n324) );
  NAND3_X1 U301 ( .A1(n322), .A2(n323), .A3(n324), .ZN(n112) );
  NOR2_X1 U302 ( .A1(n113), .A2(n118), .ZN(n326) );
  XOR2_X1 U303 ( .A(n244), .B(a[6]), .Z(n327) );
  NOR2_X1 U304 ( .A1(n113), .A2(n118), .ZN(n52) );
  BUF_X2 U305 ( .A(n227), .Z(n351) );
  NAND2_X1 U306 ( .A1(n334), .A2(n237), .ZN(n328) );
  NAND2_X1 U307 ( .A1(n334), .A2(n305), .ZN(n233) );
  BUF_X2 U308 ( .A(n238), .Z(n329) );
  CLKBUF_X1 U309 ( .A(n247), .Z(n330) );
  AOI21_X1 U310 ( .B1(n303), .B2(n336), .A(n28), .ZN(n331) );
  CLKBUF_X1 U311 ( .A(n36), .Z(n332) );
  INV_X1 U312 ( .A(n350), .ZN(n333) );
  XNOR2_X1 U313 ( .A(n245), .B(a[6]), .ZN(n236) );
  NOR2_X1 U314 ( .A1(n119), .A2(n124), .ZN(n55) );
  NOR2_X1 U315 ( .A1(n96), .A2(n95), .ZN(n20) );
  XOR2_X1 U316 ( .A(n245), .B(a[4]), .Z(n334) );
  OAI21_X1 U317 ( .B1(n306), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U318 ( .A(n294), .ZN(n38) );
  INV_X1 U319 ( .A(n39), .ZN(n37) );
  INV_X1 U320 ( .A(n30), .ZN(n28) );
  AOI21_X1 U321 ( .B1(n338), .B2(n66), .A(n63), .ZN(n61) );
  NAND2_X1 U322 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U323 ( .A(n321), .ZN(n88) );
  INV_X1 U324 ( .A(n20), .ZN(n81) );
  NAND2_X1 U325 ( .A1(n335), .A2(n301), .ZN(n3) );
  XOR2_X1 U326 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U327 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U328 ( .A(n41), .ZN(n84) );
  XOR2_X1 U329 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U330 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U331 ( .A(n55), .ZN(n87) );
  XNOR2_X1 U332 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U333 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U334 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  INV_X1 U335 ( .A(n326), .ZN(n86) );
  NOR2_X1 U336 ( .A1(n107), .A2(n112), .ZN(n46) );
  XNOR2_X1 U337 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U338 ( .A1(n337), .A2(n77), .ZN(n12) );
  OR2_X1 U339 ( .A1(n169), .A2(n157), .ZN(n116) );
  NOR2_X1 U340 ( .A1(n103), .A2(n106), .ZN(n41) );
  NAND2_X1 U341 ( .A1(n119), .A2(n124), .ZN(n56) );
  NAND2_X1 U342 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U343 ( .A(n71), .ZN(n91) );
  INV_X1 U344 ( .A(n94), .ZN(n95) );
  XOR2_X1 U345 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U346 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U347 ( .A(n67), .ZN(n90) );
  NOR2_X1 U348 ( .A1(n125), .A2(n128), .ZN(n59) );
  INV_X1 U349 ( .A(n80), .ZN(n78) );
  NAND2_X1 U350 ( .A1(n125), .A2(n128), .ZN(n60) );
  NAND2_X1 U351 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U352 ( .A1(n182), .A2(n175), .ZN(n337) );
  NAND2_X1 U353 ( .A1(n113), .A2(n118), .ZN(n53) );
  NAND2_X1 U354 ( .A1(n103), .A2(n106), .ZN(n42) );
  AND2_X1 U355 ( .A1(n351), .A2(n143), .ZN(n175) );
  OR2_X1 U356 ( .A1(n129), .A2(n132), .ZN(n338) );
  INV_X1 U357 ( .A(n14), .ZN(product[15]) );
  AND2_X1 U358 ( .A1(n351), .A2(n140), .ZN(n167) );
  OR2_X1 U359 ( .A1(n351), .A2(n241), .ZN(n201) );
  INV_X1 U360 ( .A(n136), .ZN(n152) );
  INV_X1 U361 ( .A(n139), .ZN(n160) );
  INV_X1 U362 ( .A(n290), .ZN(n101) );
  AND2_X1 U363 ( .A1(n351), .A2(n350), .ZN(n159) );
  NOR2_X1 U364 ( .A1(n133), .A2(n134), .ZN(n67) );
  NAND2_X1 U365 ( .A1(n133), .A2(n134), .ZN(n68) );
  AND2_X1 U366 ( .A1(n286), .A2(n80), .ZN(product[1]) );
  OR2_X1 U367 ( .A1(n351), .A2(n240), .ZN(n192) );
  OR2_X1 U368 ( .A1(n351), .A2(n242), .ZN(n210) );
  OR2_X1 U369 ( .A1(n351), .A2(n243), .ZN(n219) );
  AND2_X1 U370 ( .A1(n351), .A2(n146), .ZN(product[0]) );
  INV_X1 U371 ( .A(n145), .ZN(n176) );
  INV_X1 U372 ( .A(n110), .ZN(n111) );
  XNOR2_X1 U373 ( .A(n244), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U374 ( .A(n244), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U375 ( .A(n244), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U376 ( .A(n351), .B(n244), .ZN(n191) );
  INV_X1 U377 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U378 ( .A(n246), .B(a[4]), .ZN(n237) );
  NAND2_X1 U379 ( .A1(n247), .A2(n342), .ZN(n343) );
  NAND2_X1 U380 ( .A1(n341), .A2(n146), .ZN(n344) );
  NAND2_X1 U381 ( .A1(n343), .A2(n344), .ZN(n231) );
  INV_X1 U382 ( .A(n247), .ZN(n341) );
  INV_X1 U383 ( .A(n146), .ZN(n342) );
  NAND2_X1 U384 ( .A1(n182), .A2(n175), .ZN(n77) );
  CLKBUF_X1 U385 ( .A(b[7]), .Z(n345) );
  NAND2_X1 U386 ( .A1(n230), .A2(n238), .ZN(n346) );
  NAND2_X1 U387 ( .A1(n230), .A2(n329), .ZN(n347) );
  NAND2_X1 U388 ( .A1(n230), .A2(n320), .ZN(n234) );
  XNOR2_X1 U389 ( .A(n247), .B(a[2]), .ZN(n238) );
  INV_X1 U390 ( .A(n142), .ZN(n168) );
  NAND2_X1 U391 ( .A1(n98), .A2(n97), .ZN(n30) );
  OAI21_X1 U392 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  INV_X1 U393 ( .A(n65), .ZN(n63) );
  NAND2_X1 U394 ( .A1(n338), .A2(n65), .ZN(n9) );
  NOR2_X1 U395 ( .A1(n46), .A2(n41), .ZN(n39) );
  INV_X1 U396 ( .A(n46), .ZN(n85) );
  NOR2_X1 U397 ( .A1(n25), .A2(n20), .ZN(n18) );
  OAI22_X1 U398 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  NAND2_X1 U399 ( .A1(n151), .A2(n183), .ZN(n80) );
  OAI22_X1 U400 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U401 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OAI22_X1 U402 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U403 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  OAI22_X1 U404 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OAI22_X1 U405 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U406 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  NAND2_X1 U407 ( .A1(n327), .A2(n236), .ZN(n348) );
  NAND2_X1 U408 ( .A1(n228), .A2(n236), .ZN(n349) );
  XOR2_X1 U409 ( .A(n245), .B(a[6]), .Z(n350) );
  XOR2_X1 U410 ( .A(n244), .B(a[6]), .Z(n228) );
  NAND2_X1 U411 ( .A1(n228), .A2(n236), .ZN(n232) );
  INV_X1 U412 ( .A(n47), .ZN(n45) );
  OAI21_X1 U413 ( .B1(n302), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U414 ( .A1(n85), .A2(n47), .ZN(n5) );
  NAND2_X1 U415 ( .A1(n107), .A2(n112), .ZN(n47) );
  NAND2_X1 U416 ( .A1(n335), .A2(n336), .ZN(n25) );
  XNOR2_X1 U417 ( .A(n9), .B(n311), .ZN(product[5]) );
  OAI21_X1 U418 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  OAI21_X1 U419 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  XOR2_X1 U420 ( .A(n11), .B(n73), .Z(product[3]) );
  AOI21_X1 U421 ( .B1(n337), .B2(n78), .A(n75), .ZN(n73) );
  OAI22_X1 U422 ( .A1(n184), .A2(n348), .B1(n184), .B2(n333), .ZN(n136) );
  OAI22_X1 U423 ( .A1(n349), .A2(n185), .B1(n184), .B2(n333), .ZN(n94) );
  OAI22_X1 U424 ( .A1(n348), .A2(n188), .B1(n187), .B2(n333), .ZN(n155) );
  OAI22_X1 U425 ( .A1(n349), .A2(n187), .B1(n186), .B2(n333), .ZN(n154) );
  OAI22_X1 U426 ( .A1(n349), .A2(n190), .B1(n189), .B2(n333), .ZN(n157) );
  OAI22_X1 U427 ( .A1(n348), .A2(n186), .B1(n185), .B2(n333), .ZN(n153) );
  OAI22_X1 U428 ( .A1(n348), .A2(n189), .B1(n188), .B2(n333), .ZN(n156) );
  OAI22_X1 U429 ( .A1(n232), .A2(n240), .B1(n192), .B2(n236), .ZN(n148) );
  OAI22_X1 U430 ( .A1(n232), .A2(n191), .B1(n190), .B2(n236), .ZN(n158) );
  XNOR2_X1 U431 ( .A(n325), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U432 ( .A(n351), .B(n325), .ZN(n200) );
  XNOR2_X1 U433 ( .A(n325), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U434 ( .A(n325), .B(b[6]), .ZN(n194) );
  INV_X1 U435 ( .A(n245), .ZN(n241) );
  INV_X1 U436 ( .A(n70), .ZN(n69) );
  INV_X1 U437 ( .A(n77), .ZN(n75) );
  OAI22_X1 U438 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  NAND2_X2 U439 ( .A1(n231), .A2(n255), .ZN(n235) );
  AOI21_X1 U440 ( .B1(n285), .B2(n336), .A(n28), .ZN(n26) );
  OAI21_X1 U441 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  INV_X1 U442 ( .A(n331), .ZN(n24) );
  OAI21_X1 U443 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  NOR2_X1 U444 ( .A1(n326), .A2(n55), .ZN(n50) );
  INV_X1 U445 ( .A(n58), .ZN(n57) );
  NAND2_X1 U446 ( .A1(n129), .A2(n132), .ZN(n65) );
  OAI22_X1 U447 ( .A1(n292), .A2(n199), .B1(n198), .B2(n340), .ZN(n165) );
  OAI22_X1 U448 ( .A1(n328), .A2(n194), .B1(n193), .B2(n340), .ZN(n100) );
  OAI22_X1 U449 ( .A1(n292), .A2(n197), .B1(n196), .B2(n304), .ZN(n163) );
  OAI22_X1 U450 ( .A1(n193), .A2(n292), .B1(n193), .B2(n340), .ZN(n139) );
  OAI22_X1 U451 ( .A1(n328), .A2(n198), .B1(n197), .B2(n304), .ZN(n164) );
  OAI22_X1 U452 ( .A1(n328), .A2(n196), .B1(n195), .B2(n304), .ZN(n162) );
  INV_X1 U453 ( .A(n340), .ZN(n140) );
  OAI22_X1 U454 ( .A1(n233), .A2(n195), .B1(n194), .B2(n304), .ZN(n161) );
  INV_X1 U455 ( .A(n318), .ZN(n242) );
  OAI22_X1 U456 ( .A1(n233), .A2(n241), .B1(n201), .B2(n304), .ZN(n149) );
  OAI22_X1 U457 ( .A1(n233), .A2(n200), .B1(n199), .B2(n340), .ZN(n166) );
  XNOR2_X1 U458 ( .A(n293), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U459 ( .A(n318), .B(b[5]), .ZN(n204) );
  XNOR2_X1 U460 ( .A(n351), .B(n318), .ZN(n209) );
  XNOR2_X1 U461 ( .A(n246), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U462 ( .A(n330), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U463 ( .A(n316), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U464 ( .A(n330), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U465 ( .A(n351), .B(n330), .ZN(n218) );
  INV_X1 U466 ( .A(n316), .ZN(n243) );
  NAND2_X1 U467 ( .A1(n39), .A2(n18), .ZN(n16) );
  AOI21_X1 U468 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XNOR2_X1 U469 ( .A(n244), .B(n345), .ZN(n184) );
  XNOR2_X1 U470 ( .A(n325), .B(n345), .ZN(n193) );
  XNOR2_X1 U471 ( .A(n316), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U472 ( .A(n246), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U473 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U474 ( .A(n8), .B(n317), .Z(product[6]) );
  AOI21_X1 U475 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  NOR2_X1 U476 ( .A1(n135), .A2(n150), .ZN(n71) );
  NAND2_X1 U477 ( .A1(n135), .A2(n150), .ZN(n72) );
  XNOR2_X1 U478 ( .A(n293), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U479 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U480 ( .A(n325), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U481 ( .A(n316), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U482 ( .A(n244), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U483 ( .A(n318), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U484 ( .A(n325), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U485 ( .A(n330), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U486 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U487 ( .A(n245), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U488 ( .A(n293), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U489 ( .A(n316), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U490 ( .A(n332), .B(n3), .ZN(product[11]) );
  AOI21_X1 U491 ( .B1(n36), .B2(n335), .A(n303), .ZN(n31) );
  AOI21_X1 U492 ( .B1(n36), .B2(n296), .A(n24), .ZN(n22) );
  OAI21_X1 U493 ( .B1(n49), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U494 ( .A(n306), .ZN(n48) );
  OAI22_X1 U495 ( .A1(n346), .A2(n204), .B1(n203), .B2(n329), .ZN(n169) );
  OAI22_X1 U496 ( .A1(n347), .A2(n207), .B1(n206), .B2(n291), .ZN(n172) );
  OAI22_X1 U497 ( .A1(n319), .A2(n206), .B1(n205), .B2(n291), .ZN(n171) );
  OAI22_X1 U498 ( .A1(n319), .A2(n205), .B1(n204), .B2(n291), .ZN(n170) );
  OAI22_X1 U499 ( .A1(n347), .A2(n208), .B1(n207), .B2(n329), .ZN(n173) );
  OAI22_X1 U500 ( .A1(n319), .A2(n242), .B1(n210), .B2(n329), .ZN(n150) );
  OAI22_X1 U501 ( .A1(n234), .A2(n203), .B1(n202), .B2(n320), .ZN(n110) );
  OAI22_X1 U502 ( .A1(n346), .A2(n202), .B1(n202), .B2(n329), .ZN(n142) );
  INV_X1 U503 ( .A(n329), .ZN(n143) );
  OAI22_X1 U504 ( .A1(n319), .A2(n209), .B1(n208), .B2(n291), .ZN(n174) );
  INV_X2 U505 ( .A(n146), .ZN(n255) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  OR2_X1 U106 ( .A1(A[0]), .A2(B[0]), .ZN(n142) );
  AOI21_X1 U107 ( .B1(n51), .B2(n151), .A(n48), .ZN(n143) );
  CLKBUF_X1 U108 ( .A(n35), .Z(n144) );
  CLKBUF_X1 U109 ( .A(n43), .Z(n145) );
  CLKBUF_X1 U110 ( .A(n27), .Z(n146) );
  AOI21_X1 U111 ( .B1(n144), .B2(n154), .A(n32), .ZN(n147) );
  AOI21_X1 U112 ( .B1(n145), .B2(n153), .A(n40), .ZN(n148) );
  XNOR2_X1 U113 ( .A(n16), .B(n149), .ZN(SUM[15]) );
  XOR2_X1 U114 ( .A(B[15]), .B(A[15]), .Z(n149) );
  INV_X1 U115 ( .A(n42), .ZN(n40) );
  INV_X1 U116 ( .A(n34), .ZN(n32) );
  INV_X1 U117 ( .A(n66), .ZN(n64) );
  AOI21_X1 U118 ( .B1(n59), .B2(n152), .A(n56), .ZN(n54) );
  INV_X1 U119 ( .A(n58), .ZN(n56) );
  OAI21_X1 U120 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  AOI21_X1 U121 ( .B1(n51), .B2(n151), .A(n48), .ZN(n46) );
  INV_X1 U122 ( .A(n50), .ZN(n48) );
  NAND2_X1 U123 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U124 ( .A(n28), .ZN(n76) );
  NAND2_X1 U125 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U126 ( .A(n52), .ZN(n82) );
  NAND2_X1 U127 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U128 ( .A(n44), .ZN(n80) );
  NAND2_X1 U129 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U130 ( .A(n36), .ZN(n78) );
  NAND2_X1 U131 ( .A1(n152), .A2(n58), .ZN(n11) );
  NAND2_X1 U132 ( .A1(n155), .A2(n26), .ZN(n3) );
  NAND2_X1 U133 ( .A1(n154), .A2(n34), .ZN(n5) );
  NAND2_X1 U134 ( .A1(n150), .A2(n66), .ZN(n13) );
  NAND2_X1 U135 ( .A1(n151), .A2(n50), .ZN(n9) );
  NAND2_X1 U136 ( .A1(n153), .A2(n42), .ZN(n7) );
  NAND2_X1 U137 ( .A1(n86), .A2(n69), .ZN(n14) );
  XNOR2_X1 U138 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  NAND2_X1 U139 ( .A1(n156), .A2(n20), .ZN(n2) );
  NAND2_X1 U140 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U141 ( .A(n60), .ZN(n84) );
  INV_X1 U142 ( .A(n20), .ZN(n18) );
  OR2_X1 U143 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  NOR2_X1 U144 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  OR2_X1 U145 ( .A1(A[6]), .A2(B[6]), .ZN(n151) );
  OR2_X1 U146 ( .A1(A[4]), .A2(B[4]), .ZN(n152) );
  NOR2_X1 U147 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U148 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U149 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NOR2_X1 U150 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NAND2_X1 U151 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U152 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U153 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U154 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U155 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U156 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  NAND2_X1 U157 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  OR2_X1 U158 ( .A1(A[8]), .A2(B[8]), .ZN(n153) );
  OR2_X1 U159 ( .A1(A[10]), .A2(B[10]), .ZN(n154) );
  OR2_X1 U160 ( .A1(A[12]), .A2(B[12]), .ZN(n155) );
  OR2_X1 U161 ( .A1(A[14]), .A2(B[14]), .ZN(n156) );
  NAND2_X1 U162 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U163 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  NAND2_X1 U164 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U165 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  INV_X1 U166 ( .A(n26), .ZN(n24) );
  AND2_X1 U167 ( .A1(n142), .A2(n71), .ZN(SUM[0]) );
  INV_X1 U168 ( .A(n22), .ZN(n73) );
  NAND2_X1 U169 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  NOR2_X1 U170 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  XNOR2_X1 U171 ( .A(n67), .B(n13), .ZN(SUM[2]) );
  XOR2_X1 U172 ( .A(n62), .B(n12), .Z(SUM[3]) );
  XOR2_X1 U173 ( .A(n14), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U174 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  AOI21_X1 U175 ( .B1(n67), .B2(n150), .A(n64), .ZN(n62) );
  XNOR2_X1 U176 ( .A(n146), .B(n3), .ZN(SUM[12]) );
  AOI21_X1 U177 ( .B1(n43), .B2(n153), .A(n40), .ZN(n38) );
  XNOR2_X1 U178 ( .A(n145), .B(n7), .ZN(SUM[8]) );
  XOR2_X1 U179 ( .A(n147), .B(n4), .Z(SUM[11]) );
  XOR2_X1 U180 ( .A(n143), .B(n8), .Z(SUM[7]) );
  INV_X1 U181 ( .A(n68), .ZN(n86) );
  OAI21_X1 U182 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U183 ( .B1(n35), .B2(n154), .A(n32), .ZN(n30) );
  OAI21_X1 U184 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  OAI21_X1 U185 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  XNOR2_X1 U186 ( .A(n144), .B(n5), .ZN(SUM[10]) );
  XNOR2_X1 U187 ( .A(n51), .B(n9), .ZN(SUM[6]) );
  XOR2_X1 U188 ( .A(n148), .B(n6), .Z(SUM[9]) );
  OAI21_X1 U189 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  XNOR2_X1 U190 ( .A(n59), .B(n11), .ZN(SUM[4]) );
  XOR2_X1 U191 ( .A(n54), .B(n10), .Z(SUM[5]) );
  OAI21_X1 U192 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X1 U193 ( .B1(n21), .B2(n156), .A(n18), .ZN(n16) );
  NAND2_X1 U194 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  AOI21_X1 U195 ( .B1(n27), .B2(n155), .A(n24), .ZN(n22) );
endmodule


module add_layer_WIDTH16_0 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_0_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_11_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  AND2_X1 U106 ( .A1(n157), .A2(n71), .ZN(SUM[0]) );
  OAI21_X1 U107 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  CLKBUF_X1 U108 ( .A(n46), .Z(n143) );
  CLKBUF_X1 U109 ( .A(n67), .Z(n144) );
  CLKBUF_X1 U110 ( .A(n27), .Z(n145) );
  AOI21_X1 U111 ( .B1(n35), .B2(n153), .A(n32), .ZN(n146) );
  AOI21_X1 U112 ( .B1(n144), .B2(n150), .A(n64), .ZN(n147) );
  CLKBUF_X1 U113 ( .A(n54), .Z(n148) );
  XNOR2_X1 U114 ( .A(n16), .B(n149), .ZN(SUM[15]) );
  XOR2_X1 U115 ( .A(B[15]), .B(A[15]), .Z(n149) );
  OAI21_X1 U116 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  INV_X1 U117 ( .A(n34), .ZN(n32) );
  INV_X1 U118 ( .A(n42), .ZN(n40) );
  OAI21_X1 U119 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X1 U120 ( .B1(n59), .B2(n151), .A(n56), .ZN(n54) );
  INV_X1 U121 ( .A(n58), .ZN(n56) );
  AOI21_X1 U122 ( .B1(n51), .B2(n156), .A(n48), .ZN(n46) );
  INV_X1 U123 ( .A(n50), .ZN(n48) );
  AOI21_X1 U124 ( .B1(n67), .B2(n150), .A(n64), .ZN(n62) );
  INV_X1 U125 ( .A(n66), .ZN(n64) );
  NAND2_X1 U126 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U127 ( .A(n36), .ZN(n78) );
  NAND2_X1 U128 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U129 ( .A(n28), .ZN(n76) );
  NAND2_X1 U130 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U131 ( .A(n60), .ZN(n84) );
  NAND2_X1 U132 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U133 ( .A(n52), .ZN(n82) );
  NAND2_X1 U134 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U135 ( .A(n44), .ZN(n80) );
  NAND2_X1 U136 ( .A1(n154), .A2(n26), .ZN(n3) );
  NAND2_X1 U137 ( .A1(n156), .A2(n50), .ZN(n9) );
  NAND2_X1 U138 ( .A1(n153), .A2(n34), .ZN(n5) );
  NAND2_X1 U139 ( .A1(n151), .A2(n58), .ZN(n11) );
  NAND2_X1 U140 ( .A1(n152), .A2(n42), .ZN(n7) );
  XNOR2_X1 U141 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  NAND2_X1 U142 ( .A1(n155), .A2(n20), .ZN(n2) );
  XNOR2_X1 U143 ( .A(n144), .B(n13), .ZN(SUM[2]) );
  NAND2_X1 U144 ( .A1(n150), .A2(n66), .ZN(n13) );
  NAND2_X1 U145 ( .A1(n86), .A2(n69), .ZN(n14) );
  INV_X1 U146 ( .A(n68), .ZN(n86) );
  INV_X1 U147 ( .A(n20), .ZN(n18) );
  NOR2_X1 U148 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  INV_X1 U149 ( .A(n26), .ZN(n24) );
  OR2_X1 U150 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  NOR2_X1 U151 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  OR2_X1 U152 ( .A1(A[4]), .A2(B[4]), .ZN(n151) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  NOR2_X1 U154 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U155 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NOR2_X1 U156 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NAND2_X1 U157 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U158 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U159 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U160 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U161 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U162 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  NAND2_X1 U163 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  OR2_X1 U164 ( .A1(A[8]), .A2(B[8]), .ZN(n152) );
  OR2_X1 U165 ( .A1(A[10]), .A2(B[10]), .ZN(n153) );
  OR2_X1 U166 ( .A1(A[12]), .A2(B[12]), .ZN(n154) );
  OR2_X1 U167 ( .A1(A[14]), .A2(B[14]), .ZN(n155) );
  OR2_X1 U168 ( .A1(A[6]), .A2(B[6]), .ZN(n156) );
  NAND2_X1 U169 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U170 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U171 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U172 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  OR2_X1 U173 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  NAND2_X1 U174 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  XNOR2_X1 U175 ( .A(n43), .B(n7), .ZN(SUM[8]) );
  OAI21_X1 U176 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XOR2_X1 U177 ( .A(n14), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U178 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  CLKBUF_X1 U179 ( .A(n38), .Z(n158) );
  AOI21_X1 U180 ( .B1(n43), .B2(n152), .A(n40), .ZN(n38) );
  XOR2_X1 U181 ( .A(n143), .B(n8), .Z(SUM[7]) );
  XNOR2_X1 U182 ( .A(n51), .B(n9), .ZN(SUM[6]) );
  OAI21_X1 U183 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  XNOR2_X1 U184 ( .A(n59), .B(n11), .ZN(SUM[4]) );
  XOR2_X1 U185 ( .A(n148), .B(n10), .Z(SUM[5]) );
  XNOR2_X1 U186 ( .A(n35), .B(n5), .ZN(SUM[10]) );
  XOR2_X1 U187 ( .A(n147), .B(n12), .Z(SUM[3]) );
  AOI21_X1 U188 ( .B1(n35), .B2(n153), .A(n32), .ZN(n30) );
  XNOR2_X1 U189 ( .A(n145), .B(n3), .ZN(SUM[12]) );
  XOR2_X1 U190 ( .A(n158), .B(n6), .Z(SUM[9]) );
  INV_X1 U191 ( .A(n22), .ZN(n73) );
  NAND2_X1 U192 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  AOI21_X1 U193 ( .B1(n27), .B2(n154), .A(n24), .ZN(n22) );
  OAI21_X1 U194 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U195 ( .B1(n21), .B2(n155), .A(n18), .ZN(n16) );
  XOR2_X1 U196 ( .A(n146), .B(n4), .Z(SUM[11]) );
endmodule


module add_layer_WIDTH16_11 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_11_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37,
         n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70,
         n71, n73, n75, n77, n79, n81, n82, n83, n84, n140, n141, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n71), .CO(n16), .S(SUM[14]) );
  NAND2_X1 U104 ( .A1(A[2]), .A2(B[2]), .ZN(n64) );
  XNOR2_X1 U105 ( .A(B[15]), .B(A[15]), .ZN(n140) );
  OR2_X1 U106 ( .A1(A[0]), .A2(B[0]), .ZN(n141) );
  AND2_X1 U107 ( .A1(n141), .A2(n70), .ZN(SUM[0]) );
  CLKBUF_X1 U108 ( .A(n54), .Z(n143) );
  AOI21_X1 U109 ( .B1(n143), .B2(n152), .A(n51), .ZN(n144) );
  CLKBUF_X1 U110 ( .A(n41), .Z(n145) );
  CLKBUF_X1 U111 ( .A(n57), .Z(n146) );
  CLKBUF_X1 U112 ( .A(n30), .Z(n147) );
  AOI21_X1 U113 ( .B1(n147), .B2(n153), .A(n27), .ZN(n148) );
  XNOR2_X1 U114 ( .A(n16), .B(n140), .ZN(SUM[15]) );
  NOR2_X1 U115 ( .A1(A[3]), .A2(B[3]), .ZN(n149) );
  CLKBUF_X1 U116 ( .A(n38), .Z(n150) );
  OR2_X1 U117 ( .A1(A[5]), .A2(B[5]), .ZN(n152) );
  INV_X1 U118 ( .A(n66), .ZN(n65) );
  INV_X1 U119 ( .A(n29), .ZN(n27) );
  AOI21_X1 U120 ( .B1(n54), .B2(n152), .A(n51), .ZN(n49) );
  INV_X1 U121 ( .A(n53), .ZN(n51) );
  AOI21_X1 U122 ( .B1(n58), .B2(n66), .A(n59), .ZN(n57) );
  OAI21_X1 U123 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  AOI21_X1 U124 ( .B1(n46), .B2(n155), .A(n43), .ZN(n41) );
  INV_X1 U125 ( .A(n45), .ZN(n43) );
  NAND2_X1 U126 ( .A1(n73), .A2(n24), .ZN(n3) );
  INV_X1 U127 ( .A(n23), .ZN(n73) );
  NAND2_X1 U128 ( .A1(n153), .A2(n29), .ZN(n4) );
  NAND2_X1 U129 ( .A1(n154), .A2(n21), .ZN(n2) );
  NAND2_X1 U130 ( .A1(n77), .A2(n40), .ZN(n7) );
  INV_X1 U131 ( .A(n39), .ZN(n77) );
  NAND2_X1 U132 ( .A1(n75), .A2(n32), .ZN(n5) );
  INV_X1 U133 ( .A(n31), .ZN(n75) );
  XOR2_X1 U134 ( .A(n65), .B(n13), .Z(SUM[2]) );
  NAND2_X1 U135 ( .A1(n83), .A2(n64), .ZN(n13) );
  INV_X1 U136 ( .A(n63), .ZN(n83) );
  XOR2_X1 U137 ( .A(n14), .B(n70), .Z(SUM[1]) );
  NAND2_X1 U138 ( .A1(n84), .A2(n68), .ZN(n14) );
  XOR2_X1 U139 ( .A(n146), .B(n11), .Z(SUM[4]) );
  NAND2_X1 U140 ( .A1(n81), .A2(n56), .ZN(n11) );
  INV_X1 U141 ( .A(n55), .ZN(n81) );
  XOR2_X1 U142 ( .A(n144), .B(n9), .Z(SUM[6]) );
  NAND2_X1 U143 ( .A1(n79), .A2(n48), .ZN(n9) );
  INV_X1 U144 ( .A(n47), .ZN(n79) );
  NAND2_X1 U145 ( .A1(n152), .A2(n53), .ZN(n10) );
  NAND2_X1 U146 ( .A1(n151), .A2(n37), .ZN(n6) );
  NAND2_X1 U147 ( .A1(n155), .A2(n45), .ZN(n8) );
  XNOR2_X1 U148 ( .A(n62), .B(n12), .ZN(SUM[3]) );
  NAND2_X1 U149 ( .A1(n82), .A2(n61), .ZN(n12) );
  OAI21_X1 U150 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  INV_X1 U151 ( .A(n37), .ZN(n35) );
  NOR2_X1 U152 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NAND2_X1 U153 ( .A1(A[0]), .A2(B[0]), .ZN(n70) );
  NOR2_X1 U154 ( .A1(A[1]), .A2(B[1]), .ZN(n67) );
  NOR2_X1 U155 ( .A1(A[6]), .A2(B[6]), .ZN(n47) );
  INV_X1 U156 ( .A(n21), .ZN(n19) );
  OR2_X1 U157 ( .A1(A[9]), .A2(B[9]), .ZN(n151) );
  NOR2_X1 U158 ( .A1(A[8]), .A2(B[8]), .ZN(n39) );
  NOR2_X1 U159 ( .A1(A[4]), .A2(B[4]), .ZN(n55) );
  NOR2_X1 U160 ( .A1(A[12]), .A2(B[12]), .ZN(n23) );
  NOR2_X1 U161 ( .A1(A[10]), .A2(B[10]), .ZN(n31) );
  NAND2_X1 U162 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U164 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U165 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U166 ( .A1(A[13]), .A2(B[13]), .ZN(n21) );
  NAND2_X1 U167 ( .A1(A[6]), .A2(B[6]), .ZN(n48) );
  OR2_X1 U168 ( .A1(A[11]), .A2(B[11]), .ZN(n153) );
  OR2_X1 U169 ( .A1(A[13]), .A2(B[13]), .ZN(n154) );
  OR2_X1 U170 ( .A1(A[7]), .A2(B[7]), .ZN(n155) );
  NAND2_X1 U171 ( .A1(A[8]), .A2(B[8]), .ZN(n40) );
  NAND2_X1 U172 ( .A1(A[4]), .A2(B[4]), .ZN(n56) );
  NAND2_X1 U173 ( .A1(A[12]), .A2(B[12]), .ZN(n24) );
  NAND2_X1 U174 ( .A1(A[10]), .A2(B[10]), .ZN(n32) );
  NOR2_X2 U175 ( .A1(A[2]), .A2(B[2]), .ZN(n63) );
  AOI21_X1 U176 ( .B1(n150), .B2(n151), .A(n35), .ZN(n156) );
  AOI21_X1 U177 ( .B1(n38), .B2(n151), .A(n35), .ZN(n33) );
  XNOR2_X1 U178 ( .A(n150), .B(n6), .ZN(SUM[9]) );
  XOR2_X1 U179 ( .A(n156), .B(n5), .Z(SUM[10]) );
  XOR2_X1 U180 ( .A(n145), .B(n7), .Z(SUM[8]) );
  INV_X1 U181 ( .A(n67), .ZN(n84) );
  OAI21_X1 U182 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U183 ( .B1(n67), .B2(n70), .A(n68), .ZN(n66) );
  XNOR2_X1 U184 ( .A(n147), .B(n4), .ZN(SUM[11]) );
  XNOR2_X1 U185 ( .A(n46), .B(n8), .ZN(SUM[7]) );
  AOI21_X1 U186 ( .B1(n30), .B2(n153), .A(n27), .ZN(n25) );
  OAI21_X1 U187 ( .B1(n33), .B2(n31), .A(n32), .ZN(n30) );
  XNOR2_X1 U188 ( .A(n143), .B(n10), .ZN(SUM[5]) );
  NAND2_X1 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  OAI21_X1 U190 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  INV_X1 U191 ( .A(n17), .ZN(n71) );
  INV_X1 U192 ( .A(n149), .ZN(n82) );
  NOR2_X1 U193 ( .A1(n63), .A2(n149), .ZN(n58) );
  OAI21_X1 U194 ( .B1(n60), .B2(n64), .A(n61), .ZN(n59) );
  NAND2_X1 U195 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  XNOR2_X1 U196 ( .A(n22), .B(n2), .ZN(SUM[13]) );
  AOI21_X1 U197 ( .B1(n22), .B2(n154), .A(n19), .ZN(n17) );
  OAI21_X1 U198 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
  XOR2_X1 U199 ( .A(n148), .B(n3), .Z(SUM[12]) );
endmodule


module add_layer_WIDTH16_4 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_4_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_0 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_4 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_0 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_0 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_11 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_0 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_0 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0 \genblk1[0].mult  ( .clk(clk), .ia(
        {\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15 \genblk1[1].mult  ( .clk(clk), 
        .ia({\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14 \genblk1[2].mult  ( .clk(clk), 
        .ia({\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13 \genblk1[3].mult  ( .clk(clk), 
        .ia({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_0 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n33, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86,
         n87, n88, n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n142, n143, n145, n146, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n227, n228, n229, n230, n231, n232, n233, n235,
         n236, n237, n238, n240, n241, n242, n243, n244, n245, n246, n247,
         n255, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n335, n336, n337, n338, n339,
         n340, n341, n342, n343;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n317), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n111), .B(n156), .CI(n162), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n170), .B(n177), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n166), .B(n149), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  CLKBUF_X1 U249 ( .A(n342), .Z(n285) );
  BUF_X1 U250 ( .A(n245), .Z(n303) );
  OR2_X1 U251 ( .A1(n183), .A2(n151), .ZN(n286) );
  BUF_X2 U252 ( .A(n238), .Z(n335) );
  CLKBUF_X1 U253 ( .A(n46), .Z(n287) );
  CLKBUF_X1 U254 ( .A(n203), .Z(n288) );
  INV_X1 U255 ( .A(n45), .ZN(n289) );
  INV_X1 U256 ( .A(n240), .ZN(n290) );
  CLKBUF_X1 U257 ( .A(n245), .Z(n291) );
  BUF_X1 U258 ( .A(n237), .Z(n339) );
  BUF_X1 U259 ( .A(n237), .Z(n340) );
  CLKBUF_X1 U260 ( .A(n336), .Z(n292) );
  BUF_X2 U261 ( .A(n246), .Z(n336) );
  NOR2_X1 U262 ( .A1(n25), .A2(n20), .ZN(n293) );
  NAND2_X1 U263 ( .A1(n231), .A2(n255), .ZN(n294) );
  OAI21_X2 U264 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  XNOR2_X1 U265 ( .A(n336), .B(b[7]), .ZN(n295) );
  XNOR2_X1 U266 ( .A(n336), .B(b[7]), .ZN(n296) );
  XNOR2_X1 U267 ( .A(n247), .B(a[2]), .ZN(n297) );
  CLKBUF_X1 U268 ( .A(n33), .Z(n298) );
  XOR2_X1 U269 ( .A(n244), .B(a[6]), .Z(n299) );
  XOR2_X1 U270 ( .A(n244), .B(a[6]), .Z(n300) );
  AOI21_X1 U271 ( .B1(n58), .B2(n50), .A(n51), .ZN(n301) );
  NAND2_X1 U272 ( .A1(n229), .A2(n237), .ZN(n302) );
  NAND2_X1 U273 ( .A1(n229), .A2(n237), .ZN(n233) );
  NOR2_X2 U274 ( .A1(n119), .A2(n124), .ZN(n55) );
  OAI21_X1 U275 ( .B1(n342), .B2(n37), .A(n38), .ZN(n304) );
  OAI21_X1 U276 ( .B1(n37), .B2(n285), .A(n38), .ZN(n305) );
  OAI21_X1 U277 ( .B1(n342), .B2(n37), .A(n38), .ZN(n36) );
  XNOR2_X1 U278 ( .A(n115), .B(n306), .ZN(n113) );
  XNOR2_X1 U279 ( .A(n120), .B(n117), .ZN(n306) );
  BUF_X2 U280 ( .A(n247), .Z(n307) );
  CLKBUF_X1 U281 ( .A(n56), .Z(n308) );
  BUF_X2 U282 ( .A(n227), .Z(n343) );
  NAND2_X1 U283 ( .A1(n297), .A2(n230), .ZN(n309) );
  BUF_X2 U284 ( .A(n338), .Z(n310) );
  NAND2_X1 U285 ( .A1(n245), .A2(n312), .ZN(n313) );
  NAND2_X1 U286 ( .A1(n311), .A2(a[4]), .ZN(n314) );
  NAND2_X1 U287 ( .A1(n313), .A2(n314), .ZN(n229) );
  INV_X1 U288 ( .A(n245), .ZN(n311) );
  INV_X1 U289 ( .A(a[4]), .ZN(n312) );
  OAI21_X1 U290 ( .B1(n41), .B2(n47), .A(n42), .ZN(n315) );
  NOR2_X2 U291 ( .A1(n103), .A2(n106), .ZN(n41) );
  AOI21_X1 U292 ( .B1(n298), .B2(n330), .A(n28), .ZN(n316) );
  OAI22_X1 U293 ( .A1(n309), .A2(n203), .B1(n296), .B2(n335), .ZN(n317) );
  NAND2_X1 U294 ( .A1(n115), .A2(n120), .ZN(n318) );
  NAND2_X1 U295 ( .A1(n115), .A2(n117), .ZN(n319) );
  NAND2_X1 U296 ( .A1(n120), .A2(n117), .ZN(n320) );
  NAND3_X1 U297 ( .A1(n318), .A2(n319), .A3(n320), .ZN(n112) );
  BUF_X1 U298 ( .A(n236), .Z(n321) );
  NOR2_X1 U299 ( .A1(n327), .A2(n55), .ZN(n322) );
  CLKBUF_X1 U300 ( .A(n327), .Z(n323) );
  AOI21_X1 U301 ( .B1(n333), .B2(n66), .A(n63), .ZN(n324) );
  AOI21_X1 U302 ( .B1(n333), .B2(n66), .A(n63), .ZN(n325) );
  AOI21_X1 U303 ( .B1(n333), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X1 U304 ( .B1(n59), .B2(n61), .A(n60), .ZN(n326) );
  NOR2_X1 U305 ( .A1(n118), .A2(n113), .ZN(n327) );
  NAND2_X1 U306 ( .A1(n299), .A2(n236), .ZN(n328) );
  NAND2_X1 U307 ( .A1(n300), .A2(n338), .ZN(n329) );
  INV_X1 U308 ( .A(n39), .ZN(n37) );
  INV_X1 U309 ( .A(n315), .ZN(n38) );
  NAND2_X1 U310 ( .A1(n85), .A2(n289), .ZN(n5) );
  INV_X1 U311 ( .A(n287), .ZN(n85) );
  INV_X1 U312 ( .A(n47), .ZN(n45) );
  INV_X1 U313 ( .A(n25), .ZN(n23) );
  INV_X1 U314 ( .A(n316), .ZN(n24) );
  AOI21_X1 U315 ( .B1(n332), .B2(n78), .A(n75), .ZN(n73) );
  NOR2_X1 U316 ( .A1(n107), .A2(n112), .ZN(n46) );
  NAND2_X1 U317 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U318 ( .A(n71), .ZN(n91) );
  NAND2_X1 U319 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U320 ( .A(n59), .ZN(n88) );
  NAND2_X1 U321 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U322 ( .A(n20), .ZN(n81) );
  NAND2_X1 U323 ( .A1(n330), .A2(n30), .ZN(n2) );
  AOI21_X1 U324 ( .B1(n33), .B2(n330), .A(n28), .ZN(n26) );
  INV_X1 U325 ( .A(n30), .ZN(n28) );
  NAND2_X1 U326 ( .A1(n331), .A2(n35), .ZN(n3) );
  XOR2_X1 U327 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U328 ( .A1(n87), .A2(n308), .ZN(n7) );
  INV_X1 U329 ( .A(n55), .ZN(n87) );
  XOR2_X1 U330 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U331 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U332 ( .A(n80), .ZN(n78) );
  XNOR2_X1 U333 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U334 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U335 ( .B1(n57), .B2(n55), .A(n308), .ZN(n54) );
  INV_X1 U336 ( .A(n323), .ZN(n86) );
  XNOR2_X1 U337 ( .A(n9), .B(n66), .ZN(product[5]) );
  NAND2_X1 U338 ( .A1(n333), .A2(n65), .ZN(n9) );
  INV_X1 U339 ( .A(n35), .ZN(n33) );
  INV_X1 U340 ( .A(n70), .ZN(n69) );
  NOR2_X1 U341 ( .A1(n327), .A2(n55), .ZN(n50) );
  XNOR2_X1 U342 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U343 ( .A1(n332), .A2(n77), .ZN(n12) );
  XOR2_X1 U344 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U345 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U346 ( .A(n67), .ZN(n90) );
  NOR2_X1 U347 ( .A1(n113), .A2(n118), .ZN(n52) );
  XNOR2_X1 U348 ( .A(n169), .B(n157), .ZN(n117) );
  INV_X1 U349 ( .A(n94), .ZN(n95) );
  OR2_X1 U350 ( .A1(n98), .A2(n97), .ZN(n330) );
  OR2_X1 U351 ( .A1(n169), .A2(n157), .ZN(n116) );
  NOR2_X1 U352 ( .A1(n96), .A2(n95), .ZN(n20) );
  NOR2_X1 U353 ( .A1(n133), .A2(n134), .ZN(n67) );
  NAND2_X1 U354 ( .A1(n119), .A2(n124), .ZN(n56) );
  NOR2_X1 U355 ( .A1(n125), .A2(n128), .ZN(n59) );
  NAND2_X1 U356 ( .A1(n113), .A2(n118), .ZN(n53) );
  NOR2_X1 U357 ( .A1(n135), .A2(n150), .ZN(n71) );
  OR2_X1 U358 ( .A1(n99), .A2(n102), .ZN(n331) );
  OR2_X1 U359 ( .A1(n182), .A2(n175), .ZN(n332) );
  OR2_X1 U360 ( .A1(n129), .A2(n132), .ZN(n333) );
  NAND2_X1 U361 ( .A1(n129), .A2(n132), .ZN(n65) );
  NAND2_X1 U362 ( .A1(n125), .A2(n128), .ZN(n60) );
  NAND2_X1 U363 ( .A1(n133), .A2(n134), .ZN(n68) );
  NAND2_X1 U364 ( .A1(n96), .A2(n95), .ZN(n21) );
  NAND2_X1 U365 ( .A1(n103), .A2(n106), .ZN(n42) );
  AND2_X1 U366 ( .A1(n343), .A2(n143), .ZN(n175) );
  INV_X1 U367 ( .A(n14), .ZN(product[15]) );
  AND2_X1 U368 ( .A1(n286), .A2(n80), .ZN(product[1]) );
  OR2_X1 U369 ( .A1(n343), .A2(n242), .ZN(n210) );
  OR2_X1 U370 ( .A1(n343), .A2(n243), .ZN(n219) );
  AND2_X1 U371 ( .A1(n343), .A2(n140), .ZN(n167) );
  INV_X1 U372 ( .A(n139), .ZN(n160) );
  INV_X1 U373 ( .A(n100), .ZN(n101) );
  AND2_X1 U374 ( .A1(n343), .A2(n137), .ZN(n159) );
  INV_X1 U375 ( .A(n145), .ZN(n176) );
  INV_X1 U376 ( .A(n136), .ZN(n152) );
  OR2_X1 U377 ( .A1(n343), .A2(n240), .ZN(n192) );
  OR2_X1 U378 ( .A1(n343), .A2(n241), .ZN(n201) );
  NAND2_X1 U379 ( .A1(n231), .A2(n255), .ZN(n235) );
  INV_X1 U380 ( .A(n146), .ZN(n255) );
  NAND2_X1 U381 ( .A1(n228), .A2(n236), .ZN(n232) );
  AND2_X1 U382 ( .A1(n343), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U383 ( .A(n247), .B(a[2]), .ZN(n238) );
  XNOR2_X1 U384 ( .A(n245), .B(a[6]), .ZN(n338) );
  OAI22_X1 U385 ( .A1(n294), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U386 ( .A1(n294), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U387 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U388 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OAI22_X1 U389 ( .A1(n294), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U390 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  NAND2_X1 U391 ( .A1(n230), .A2(n297), .ZN(n337) );
  INV_X1 U392 ( .A(n41), .ZN(n84) );
  NOR2_X1 U393 ( .A1(n46), .A2(n41), .ZN(n39) );
  OAI21_X1 U394 ( .B1(n41), .B2(n47), .A(n42), .ZN(n40) );
  XNOR2_X1 U395 ( .A(n245), .B(a[6]), .ZN(n236) );
  XNOR2_X1 U396 ( .A(n343), .B(n244), .ZN(n191) );
  XOR2_X1 U397 ( .A(n244), .B(a[6]), .Z(n228) );
  INV_X1 U398 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U399 ( .A(n290), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U400 ( .A(n290), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U401 ( .A(n290), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U402 ( .A(n244), .B(b[3]), .ZN(n188) );
  INV_X1 U403 ( .A(n65), .ZN(n63) );
  XNOR2_X1 U404 ( .A(n246), .B(a[4]), .ZN(n237) );
  XNOR2_X1 U405 ( .A(n290), .B(b[6]), .ZN(n185) );
  CLKBUF_X1 U406 ( .A(n247), .Z(n341) );
  AOI21_X1 U407 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  OAI21_X1 U408 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U409 ( .A1(n98), .A2(n97), .ZN(n30) );
  XOR2_X1 U410 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U411 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  NAND2_X1 U412 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U413 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OAI22_X1 U414 ( .A1(n294), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  XNOR2_X1 U415 ( .A(n244), .B(b[2]), .ZN(n189) );
  INV_X1 U416 ( .A(n110), .ZN(n111) );
  NAND2_X1 U417 ( .A1(n107), .A2(n112), .ZN(n47) );
  NAND2_X1 U418 ( .A1(n135), .A2(n150), .ZN(n72) );
  OAI22_X1 U419 ( .A1(n211), .A2(n294), .B1(n211), .B2(n255), .ZN(n145) );
  OAI21_X1 U420 ( .B1(n59), .B2(n324), .A(n60), .ZN(n58) );
  INV_X1 U421 ( .A(n77), .ZN(n75) );
  AOI21_X1 U422 ( .B1(n322), .B2(n326), .A(n51), .ZN(n342) );
  NAND2_X1 U423 ( .A1(n99), .A2(n102), .ZN(n35) );
  OAI21_X1 U424 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  INV_X1 U425 ( .A(n142), .ZN(n168) );
  XOR2_X1 U426 ( .A(n22), .B(n1), .Z(product[13]) );
  OAI22_X1 U427 ( .A1(n184), .A2(n329), .B1(n184), .B2(n310), .ZN(n136) );
  OAI22_X1 U428 ( .A1(n328), .A2(n185), .B1(n184), .B2(n310), .ZN(n94) );
  OAI22_X1 U429 ( .A1(n232), .A2(n188), .B1(n187), .B2(n310), .ZN(n155) );
  OAI22_X1 U430 ( .A1(n329), .A2(n187), .B1(n186), .B2(n310), .ZN(n154) );
  INV_X1 U431 ( .A(n338), .ZN(n137) );
  OAI22_X1 U432 ( .A1(n328), .A2(n186), .B1(n185), .B2(n310), .ZN(n153) );
  OAI22_X1 U433 ( .A1(n232), .A2(n190), .B1(n189), .B2(n338), .ZN(n157) );
  OAI22_X1 U434 ( .A1(n329), .A2(n189), .B1(n188), .B2(n338), .ZN(n156) );
  XNOR2_X1 U435 ( .A(n303), .B(b[2]), .ZN(n198) );
  OAI22_X1 U436 ( .A1(n232), .A2(n240), .B1(n192), .B2(n321), .ZN(n148) );
  OAI22_X1 U437 ( .A1(n328), .A2(n191), .B1(n190), .B2(n321), .ZN(n158) );
  XNOR2_X1 U438 ( .A(n303), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U439 ( .A(n343), .B(n303), .ZN(n200) );
  XNOR2_X1 U440 ( .A(n303), .B(b[4]), .ZN(n196) );
  INV_X1 U441 ( .A(n245), .ZN(n241) );
  XNOR2_X1 U442 ( .A(n303), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U443 ( .A(n291), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U444 ( .A(n291), .B(b[6]), .ZN(n194) );
  NOR2_X1 U445 ( .A1(n25), .A2(n20), .ZN(n18) );
  NAND2_X1 U446 ( .A1(n331), .A2(n330), .ZN(n25) );
  NAND2_X1 U447 ( .A1(n39), .A2(n293), .ZN(n16) );
  XOR2_X1 U448 ( .A(n31), .B(n2), .Z(product[12]) );
  INV_X1 U449 ( .A(n326), .ZN(n57) );
  OAI22_X1 U450 ( .A1(n302), .A2(n199), .B1(n198), .B2(n339), .ZN(n165) );
  OAI22_X1 U451 ( .A1(n233), .A2(n197), .B1(n196), .B2(n340), .ZN(n163) );
  OAI22_X1 U452 ( .A1(n302), .A2(n198), .B1(n197), .B2(n339), .ZN(n164) );
  OAI22_X1 U453 ( .A1(n302), .A2(n194), .B1(n193), .B2(n340), .ZN(n100) );
  OAI22_X1 U454 ( .A1(n302), .A2(n196), .B1(n195), .B2(n339), .ZN(n162) );
  INV_X1 U455 ( .A(n340), .ZN(n140) );
  OAI22_X1 U456 ( .A1(n193), .A2(n302), .B1(n193), .B2(n339), .ZN(n139) );
  OAI22_X1 U457 ( .A1(n233), .A2(n241), .B1(n201), .B2(n340), .ZN(n149) );
  OAI22_X1 U458 ( .A1(n233), .A2(n195), .B1(n194), .B2(n339), .ZN(n161) );
  OAI22_X1 U459 ( .A1(n233), .A2(n200), .B1(n199), .B2(n340), .ZN(n166) );
  XNOR2_X1 U460 ( .A(n336), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U461 ( .A(n292), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U462 ( .A(n336), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U463 ( .A(n336), .B(b[5]), .ZN(n204) );
  INV_X1 U464 ( .A(n292), .ZN(n242) );
  XNOR2_X1 U465 ( .A(n336), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U466 ( .A(n343), .B(n336), .ZN(n209) );
  XNOR2_X1 U467 ( .A(n336), .B(b[7]), .ZN(n202) );
  XOR2_X1 U468 ( .A(n246), .B(a[2]), .Z(n230) );
  XNOR2_X1 U469 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U470 ( .A(n8), .B(n325), .Z(product[6]) );
  AOI21_X1 U471 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  NAND2_X1 U472 ( .A1(n183), .A2(n151), .ZN(n80) );
  XNOR2_X1 U473 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U474 ( .A(n291), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U475 ( .A(n336), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U476 ( .A(n305), .B(n3), .ZN(product[11]) );
  AOI21_X1 U477 ( .B1(n304), .B2(n331), .A(n298), .ZN(n31) );
  AOI21_X1 U478 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U479 ( .B1(n301), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U480 ( .A(n301), .ZN(n48) );
  OAI22_X1 U481 ( .A1(n337), .A2(n204), .B1(n288), .B2(n335), .ZN(n169) );
  OAI22_X1 U482 ( .A1(n337), .A2(n207), .B1(n206), .B2(n335), .ZN(n172) );
  OAI22_X1 U483 ( .A1(n337), .A2(n206), .B1(n205), .B2(n335), .ZN(n171) );
  OAI22_X1 U484 ( .A1(n337), .A2(n205), .B1(n204), .B2(n335), .ZN(n170) );
  OAI22_X1 U485 ( .A1(n337), .A2(n208), .B1(n207), .B2(n335), .ZN(n173) );
  OAI22_X1 U486 ( .A1(n337), .A2(n242), .B1(n210), .B2(n335), .ZN(n150) );
  OAI22_X1 U487 ( .A1(n309), .A2(n203), .B1(n296), .B2(n335), .ZN(n110) );
  XNOR2_X1 U488 ( .A(n341), .B(b[5]), .ZN(n213) );
  OAI22_X1 U489 ( .A1(n295), .A2(n309), .B1(n202), .B2(n335), .ZN(n142) );
  XNOR2_X1 U490 ( .A(n307), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U491 ( .A(n341), .B(b[4]), .ZN(n214) );
  INV_X1 U492 ( .A(n335), .ZN(n143) );
  OAI22_X1 U493 ( .A1(n309), .A2(n209), .B1(n208), .B2(n335), .ZN(n174) );
  XNOR2_X1 U494 ( .A(n307), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U495 ( .A(n343), .B(n341), .ZN(n218) );
  XNOR2_X1 U496 ( .A(n307), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U497 ( .A(n307), .B(b[2]), .ZN(n216) );
  INV_X1 U498 ( .A(n307), .ZN(n243) );
  XNOR2_X1 U499 ( .A(n307), .B(b[1]), .ZN(n217) );
  XOR2_X1 U500 ( .A(n247), .B(n146), .Z(n231) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n33, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n66, n67, n68,
         n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n87, n88,
         n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n139,
         n140, n142, n143, n145, n146, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n227, n229, n230, n231, n232, n233, n234, n235, n237, n238, n240,
         n241, n242, n243, n244, n245, n246, n247, n255, n285, n286, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n168), .CI(n334), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n156), .B(n162), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n170), .B(n164), .CI(n177), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n148), .B(n158), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  OAI21_X1 U249 ( .B1(n41), .B2(n47), .A(n42), .ZN(n285) );
  BUF_X2 U250 ( .A(n247), .Z(n343) );
  OR2_X1 U251 ( .A1(n99), .A2(n102), .ZN(n341) );
  AND2_X1 U252 ( .A1(n129), .A2(n132), .ZN(n286) );
  AND2_X1 U253 ( .A1(n338), .A2(n80), .ZN(product[1]) );
  INV_X1 U254 ( .A(n286), .ZN(n288) );
  INV_X1 U255 ( .A(n88), .ZN(n289) );
  NOR2_X1 U256 ( .A1(n125), .A2(n128), .ZN(n59) );
  CLKBUF_X1 U257 ( .A(n66), .Z(n290) );
  OAI21_X1 U258 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  CLKBUF_X1 U259 ( .A(n350), .Z(n291) );
  INV_X1 U260 ( .A(n87), .ZN(n292) );
  NAND2_X1 U261 ( .A1(n328), .A2(n329), .ZN(n293) );
  CLKBUF_X1 U262 ( .A(n56), .Z(n294) );
  CLKBUF_X1 U263 ( .A(n343), .Z(n295) );
  CLKBUF_X1 U264 ( .A(n47), .Z(n296) );
  CLKBUF_X1 U265 ( .A(n232), .Z(n346) );
  INV_X1 U266 ( .A(n140), .ZN(n297) );
  XOR2_X1 U267 ( .A(n241), .B(b[2]), .Z(n198) );
  NAND2_X1 U268 ( .A1(n231), .A2(n255), .ZN(n298) );
  BUF_X1 U269 ( .A(n238), .Z(n299) );
  CLKBUF_X1 U270 ( .A(n349), .Z(n300) );
  BUF_X2 U271 ( .A(n349), .Z(n301) );
  BUF_X1 U272 ( .A(n246), .Z(n349) );
  CLKBUF_X1 U273 ( .A(n73), .Z(n302) );
  CLKBUF_X1 U274 ( .A(n245), .Z(n303) );
  CLKBUF_X1 U275 ( .A(n151), .Z(n304) );
  OAI21_X1 U276 ( .B1(n335), .B2(n56), .A(n53), .ZN(n305) );
  XNOR2_X1 U277 ( .A(n316), .B(b[7]), .ZN(n306) );
  CLKBUF_X1 U278 ( .A(n246), .Z(n307) );
  XNOR2_X1 U279 ( .A(n247), .B(a[2]), .ZN(n308) );
  CLKBUF_X1 U280 ( .A(n245), .Z(n309) );
  XNOR2_X2 U281 ( .A(n307), .B(a[4]), .ZN(n350) );
  INV_X1 U282 ( .A(n240), .ZN(n310) );
  CLKBUF_X1 U283 ( .A(n234), .Z(n315) );
  OR2_X2 U284 ( .A1(n312), .A2(n311), .ZN(n232) );
  XNOR2_X1 U285 ( .A(n244), .B(a[6]), .ZN(n311) );
  XOR2_X1 U286 ( .A(n245), .B(a[6]), .Z(n312) );
  XNOR2_X1 U287 ( .A(n122), .B(n313), .ZN(n115) );
  XNOR2_X1 U288 ( .A(n163), .B(n176), .ZN(n313) );
  CLKBUF_X1 U289 ( .A(n246), .Z(n316) );
  CLKBUF_X1 U290 ( .A(n245), .Z(n314) );
  CLKBUF_X1 U291 ( .A(n33), .Z(n317) );
  NAND2_X1 U292 ( .A1(n229), .A2(n237), .ZN(n318) );
  NAND2_X1 U293 ( .A1(n293), .A2(n237), .ZN(n319) );
  NAND2_X1 U294 ( .A1(n293), .A2(n237), .ZN(n233) );
  NAND2_X1 U295 ( .A1(n122), .A2(n163), .ZN(n320) );
  NAND2_X1 U296 ( .A1(n122), .A2(n176), .ZN(n321) );
  NAND2_X1 U297 ( .A1(n163), .A2(n176), .ZN(n322) );
  NAND3_X1 U298 ( .A1(n320), .A2(n321), .A3(n322), .ZN(n114) );
  XNOR2_X1 U299 ( .A(n115), .B(n324), .ZN(n323) );
  XNOR2_X1 U300 ( .A(n115), .B(n324), .ZN(n113) );
  XNOR2_X1 U301 ( .A(n120), .B(n117), .ZN(n324) );
  AOI21_X1 U302 ( .B1(n342), .B2(n66), .A(n286), .ZN(n325) );
  NAND2_X1 U303 ( .A1(n245), .A2(n327), .ZN(n328) );
  NAND2_X1 U304 ( .A1(n326), .A2(a[4]), .ZN(n329) );
  NAND2_X1 U305 ( .A1(n328), .A2(n329), .ZN(n229) );
  INV_X1 U306 ( .A(n245), .ZN(n326) );
  INV_X1 U307 ( .A(a[4]), .ZN(n327) );
  AOI21_X1 U308 ( .B1(n342), .B2(n66), .A(n286), .ZN(n61) );
  NAND2_X1 U309 ( .A1(n115), .A2(n120), .ZN(n330) );
  NAND2_X1 U310 ( .A1(n115), .A2(n117), .ZN(n331) );
  NAND2_X1 U311 ( .A1(n120), .A2(n117), .ZN(n332) );
  NAND3_X1 U312 ( .A1(n330), .A2(n331), .A3(n332), .ZN(n112) );
  OAI21_X2 U313 ( .B1(n49), .B2(n37), .A(n38), .ZN(n36) );
  AOI21_X1 U314 ( .B1(n317), .B2(n340), .A(n28), .ZN(n333) );
  OAI22_X1 U315 ( .A1(n354), .A2(n203), .B1(n306), .B2(n299), .ZN(n334) );
  NOR2_X1 U316 ( .A1(n323), .A2(n118), .ZN(n335) );
  XNOR2_X1 U317 ( .A(n245), .B(a[6]), .ZN(n336) );
  XNOR2_X1 U318 ( .A(n31), .B(n337), .ZN(product[12]) );
  AND2_X1 U319 ( .A1(n340), .A2(n30), .ZN(n337) );
  NOR2_X1 U320 ( .A1(n119), .A2(n124), .ZN(n55) );
  OR2_X1 U321 ( .A1(n98), .A2(n97), .ZN(n340) );
  INV_X1 U322 ( .A(n285), .ZN(n38) );
  INV_X1 U323 ( .A(n39), .ZN(n37) );
  XNOR2_X1 U324 ( .A(n48), .B(n5), .ZN(product[9]) );
  INV_X1 U325 ( .A(n46), .ZN(n85) );
  INV_X1 U326 ( .A(n25), .ZN(n23) );
  NOR2_X1 U327 ( .A1(n107), .A2(n112), .ZN(n46) );
  AOI21_X1 U328 ( .B1(n33), .B2(n340), .A(n28), .ZN(n26) );
  INV_X1 U329 ( .A(n30), .ZN(n28) );
  NAND2_X1 U330 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U331 ( .A(n59), .ZN(n88) );
  NAND2_X1 U332 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U333 ( .A(n20), .ZN(n81) );
  AOI21_X1 U334 ( .B1(n339), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U335 ( .A(n77), .ZN(n75) );
  NAND2_X1 U336 ( .A1(n342), .A2(n288), .ZN(n9) );
  XOR2_X1 U337 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U338 ( .A1(n87), .A2(n294), .ZN(n7) );
  INV_X1 U339 ( .A(n55), .ZN(n87) );
  XOR2_X1 U340 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U341 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U342 ( .A(n41), .ZN(n84) );
  XNOR2_X1 U343 ( .A(n54), .B(n6), .ZN(product[8]) );
  OAI21_X1 U344 ( .B1(n57), .B2(n292), .A(n294), .ZN(n54) );
  NOR2_X1 U345 ( .A1(n46), .A2(n41), .ZN(n39) );
  NOR2_X1 U346 ( .A1(n25), .A2(n20), .ZN(n18) );
  XNOR2_X1 U347 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U348 ( .A1(n339), .A2(n77), .ZN(n12) );
  OR2_X1 U349 ( .A1(n183), .A2(n304), .ZN(n338) );
  NOR2_X1 U350 ( .A1(n96), .A2(n95), .ZN(n20) );
  NAND2_X1 U351 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U352 ( .A(n71), .ZN(n91) );
  OR2_X1 U353 ( .A1(n169), .A2(n157), .ZN(n116) );
  INV_X1 U354 ( .A(n94), .ZN(n95) );
  XNOR2_X1 U355 ( .A(n169), .B(n157), .ZN(n117) );
  OR2_X1 U356 ( .A1(n182), .A2(n175), .ZN(n339) );
  XOR2_X1 U357 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U358 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U359 ( .A(n67), .ZN(n90) );
  NAND2_X1 U360 ( .A1(n119), .A2(n124), .ZN(n56) );
  NAND2_X1 U361 ( .A1(n125), .A2(n128), .ZN(n60) );
  NAND2_X1 U362 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U363 ( .A1(n132), .A2(n129), .ZN(n342) );
  INV_X1 U364 ( .A(n70), .ZN(n69) );
  AND2_X1 U365 ( .A1(n227), .A2(n143), .ZN(n175) );
  INV_X1 U366 ( .A(n14), .ZN(product[15]) );
  AND2_X1 U367 ( .A1(n227), .A2(n140), .ZN(n167) );
  OR2_X1 U368 ( .A1(n227), .A2(n243), .ZN(n219) );
  OR2_X1 U369 ( .A1(n227), .A2(n241), .ZN(n201) );
  INV_X1 U370 ( .A(n136), .ZN(n152) );
  INV_X1 U371 ( .A(n139), .ZN(n160) );
  INV_X1 U372 ( .A(n100), .ZN(n101) );
  INV_X1 U373 ( .A(n145), .ZN(n176) );
  INV_X1 U374 ( .A(n142), .ZN(n168) );
  AND2_X1 U375 ( .A1(n227), .A2(n347), .ZN(n159) );
  NOR2_X1 U376 ( .A1(n133), .A2(n134), .ZN(n67) );
  NAND2_X1 U377 ( .A1(n135), .A2(n150), .ZN(n72) );
  NAND2_X1 U378 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U379 ( .A1(n227), .A2(n240), .ZN(n192) );
  OR2_X1 U380 ( .A1(n227), .A2(n242), .ZN(n210) );
  INV_X1 U381 ( .A(n146), .ZN(n255) );
  NAND2_X1 U382 ( .A1(n231), .A2(n255), .ZN(n235) );
  AND2_X1 U383 ( .A1(n227), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U384 ( .A(n310), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U385 ( .A(n310), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U386 ( .A(n244), .B(b[2]), .ZN(n189) );
  INV_X1 U387 ( .A(n244), .ZN(n240) );
  BUF_X2 U388 ( .A(n238), .Z(n344) );
  XNOR2_X1 U389 ( .A(n247), .B(a[2]), .ZN(n238) );
  BUF_X2 U390 ( .A(n336), .Z(n345) );
  NAND2_X1 U391 ( .A1(n341), .A2(n340), .ZN(n25) );
  NAND2_X1 U392 ( .A1(n341), .A2(n35), .ZN(n3) );
  NOR2_X1 U393 ( .A1(n135), .A2(n150), .ZN(n71) );
  XOR2_X1 U394 ( .A(n314), .B(a[6]), .Z(n347) );
  NAND2_X1 U395 ( .A1(n103), .A2(n106), .ZN(n42) );
  NOR2_X2 U396 ( .A1(n103), .A2(n106), .ZN(n41) );
  AOI21_X1 U397 ( .B1(n50), .B2(n58), .A(n51), .ZN(n348) );
  AOI21_X1 U398 ( .B1(n50), .B2(n58), .A(n305), .ZN(n49) );
  INV_X1 U399 ( .A(n333), .ZN(n24) );
  OAI21_X1 U400 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U401 ( .A1(n98), .A2(n97), .ZN(n30) );
  XNOR2_X1 U402 ( .A(n310), .B(b[6]), .ZN(n185) );
  INV_X1 U403 ( .A(n80), .ZN(n78) );
  INV_X1 U404 ( .A(n296), .ZN(n45) );
  OAI21_X1 U405 ( .B1(n41), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U406 ( .A1(n85), .A2(n296), .ZN(n5) );
  NAND2_X1 U407 ( .A1(n107), .A2(n112), .ZN(n47) );
  OAI22_X1 U408 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U409 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U410 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  OAI22_X1 U411 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U412 ( .A1(n298), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OAI22_X1 U413 ( .A1(n211), .A2(n298), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U414 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OAI22_X1 U415 ( .A1(n298), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U416 ( .A1(n298), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  NAND2_X1 U417 ( .A1(n351), .A2(n53), .ZN(n6) );
  XNOR2_X1 U418 ( .A(n246), .B(a[4]), .ZN(n237) );
  XOR2_X1 U419 ( .A(n11), .B(n302), .Z(product[3]) );
  OAI21_X1 U420 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  NAND2_X1 U421 ( .A1(n182), .A2(n175), .ZN(n77) );
  OR2_X1 U422 ( .A1(n323), .A2(n118), .ZN(n351) );
  OR2_X1 U423 ( .A1(n232), .A2(n191), .ZN(n352) );
  OR2_X1 U424 ( .A1(n190), .A2(n336), .ZN(n353) );
  NAND2_X1 U425 ( .A1(n352), .A2(n353), .ZN(n158) );
  XNOR2_X1 U426 ( .A(n227), .B(n244), .ZN(n191) );
  XNOR2_X1 U427 ( .A(n244), .B(b[1]), .ZN(n190) );
  NAND2_X1 U428 ( .A1(n230), .A2(n308), .ZN(n354) );
  NAND2_X1 U429 ( .A1(n230), .A2(n308), .ZN(n234) );
  OAI21_X1 U430 ( .B1(n289), .B2(n325), .A(n60), .ZN(n355) );
  NAND2_X1 U431 ( .A1(n99), .A2(n102), .ZN(n35) );
  INV_X1 U432 ( .A(n110), .ZN(n111) );
  INV_X1 U433 ( .A(n35), .ZN(n33) );
  INV_X1 U434 ( .A(n355), .ZN(n57) );
  OAI21_X1 U435 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  XOR2_X1 U436 ( .A(n8), .B(n325), .Z(product[6]) );
  XNOR2_X1 U437 ( .A(n310), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U438 ( .A(n9), .B(n290), .ZN(product[5]) );
  OAI22_X1 U439 ( .A1(n319), .A2(n199), .B1(n198), .B2(n297), .ZN(n165) );
  OAI22_X1 U440 ( .A1(n319), .A2(n197), .B1(n196), .B2(n291), .ZN(n163) );
  OAI22_X1 U441 ( .A1(n318), .A2(n198), .B1(n197), .B2(n350), .ZN(n164) );
  OAI22_X1 U442 ( .A1(n319), .A2(n194), .B1(n193), .B2(n291), .ZN(n100) );
  OAI22_X1 U443 ( .A1(n193), .A2(n319), .B1(n193), .B2(n297), .ZN(n139) );
  OAI22_X1 U444 ( .A1(n318), .A2(n196), .B1(n195), .B2(n350), .ZN(n162) );
  OAI22_X1 U445 ( .A1(n233), .A2(n241), .B1(n201), .B2(n350), .ZN(n149) );
  OAI22_X1 U446 ( .A1(n318), .A2(n195), .B1(n194), .B2(n350), .ZN(n161) );
  INV_X1 U447 ( .A(n350), .ZN(n140) );
  OAI22_X1 U448 ( .A1(n233), .A2(n200), .B1(n199), .B2(n350), .ZN(n166) );
  XNOR2_X1 U449 ( .A(n301), .B(b[5]), .ZN(n204) );
  XNOR2_X1 U450 ( .A(n300), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U451 ( .A(n301), .B(b[2]), .ZN(n207) );
  INV_X1 U452 ( .A(n301), .ZN(n242) );
  XNOR2_X1 U453 ( .A(n316), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U454 ( .A(n316), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U455 ( .A(n227), .B(n301), .ZN(n209) );
  XNOR2_X1 U456 ( .A(n300), .B(b[1]), .ZN(n208) );
  XOR2_X1 U457 ( .A(n246), .B(a[2]), .Z(n230) );
  XOR2_X1 U458 ( .A(n22), .B(n1), .Z(product[13]) );
  NAND2_X1 U459 ( .A1(n151), .A2(n183), .ZN(n80) );
  OAI22_X1 U460 ( .A1(n184), .A2(n346), .B1(n184), .B2(n345), .ZN(n136) );
  NOR2_X1 U461 ( .A1(n52), .A2(n55), .ZN(n50) );
  OAI21_X1 U462 ( .B1(n335), .B2(n56), .A(n53), .ZN(n51) );
  NAND2_X1 U463 ( .A1(n113), .A2(n118), .ZN(n53) );
  NOR2_X1 U464 ( .A1(n113), .A2(n118), .ZN(n52) );
  OAI22_X1 U465 ( .A1(n346), .A2(n185), .B1(n184), .B2(n345), .ZN(n94) );
  OAI22_X1 U466 ( .A1(n346), .A2(n188), .B1(n187), .B2(n345), .ZN(n155) );
  OAI22_X1 U467 ( .A1(n346), .A2(n187), .B1(n186), .B2(n345), .ZN(n154) );
  OAI22_X1 U468 ( .A1(n346), .A2(n186), .B1(n185), .B2(n345), .ZN(n153) );
  OAI22_X1 U469 ( .A1(n232), .A2(n190), .B1(n189), .B2(n345), .ZN(n157) );
  OAI22_X1 U470 ( .A1(n232), .A2(n189), .B1(n188), .B2(n345), .ZN(n156) );
  OAI22_X1 U471 ( .A1(n232), .A2(n240), .B1(n192), .B2(n345), .ZN(n148) );
  XNOR2_X1 U472 ( .A(n309), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U473 ( .A(n314), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U474 ( .A(n309), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U475 ( .A(n227), .B(n314), .ZN(n200) );
  XNOR2_X1 U476 ( .A(n303), .B(b[6]), .ZN(n194) );
  INV_X1 U477 ( .A(n245), .ZN(n241) );
  XNOR2_X1 U478 ( .A(n303), .B(b[1]), .ZN(n199) );
  NAND2_X1 U479 ( .A1(n18), .A2(n39), .ZN(n16) );
  AOI21_X1 U480 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XNOR2_X1 U481 ( .A(n343), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U482 ( .A(n343), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U483 ( .A(n343), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U484 ( .A(n343), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U485 ( .A(n343), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U486 ( .A(n227), .B(n295), .ZN(n218) );
  XNOR2_X1 U487 ( .A(n343), .B(b[1]), .ZN(n217) );
  INV_X1 U488 ( .A(n343), .ZN(n243) );
  XOR2_X1 U489 ( .A(n247), .B(n146), .Z(n231) );
  XNOR2_X1 U490 ( .A(n301), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U491 ( .A(n309), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U492 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U493 ( .A(n343), .B(b[3]), .ZN(n215) );
  AOI21_X1 U494 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  XNOR2_X1 U495 ( .A(n36), .B(n3), .ZN(product[11]) );
  AOI21_X1 U496 ( .B1(n36), .B2(n341), .A(n317), .ZN(n31) );
  AOI21_X1 U497 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U498 ( .B1(n348), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U499 ( .A(n348), .ZN(n48) );
  OAI22_X1 U500 ( .A1(n315), .A2(n204), .B1(n203), .B2(n299), .ZN(n169) );
  OAI22_X1 U501 ( .A1(n354), .A2(n207), .B1(n206), .B2(n344), .ZN(n172) );
  OAI22_X1 U502 ( .A1(n354), .A2(n206), .B1(n205), .B2(n344), .ZN(n171) );
  OAI22_X1 U503 ( .A1(n354), .A2(n205), .B1(n204), .B2(n299), .ZN(n170) );
  OAI22_X1 U504 ( .A1(n315), .A2(n208), .B1(n207), .B2(n344), .ZN(n173) );
  OAI22_X1 U505 ( .A1(n315), .A2(n242), .B1(n210), .B2(n299), .ZN(n150) );
  OAI22_X1 U506 ( .A1(n354), .A2(n203), .B1(n202), .B2(n299), .ZN(n110) );
  OAI22_X1 U507 ( .A1(n234), .A2(n306), .B1(n202), .B2(n238), .ZN(n142) );
  INV_X1 U508 ( .A(n344), .ZN(n143) );
  OAI22_X1 U509 ( .A1(n234), .A2(n209), .B1(n208), .B2(n344), .ZN(n174) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n35, n36,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n87, n88,
         n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n139,
         n140, n142, n143, n145, n146, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n240, n241, n242, n243, n244, n245, n246, n247, n255, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n297), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n162), .B(n156), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n177), .B(n170), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n148), .B(n158), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  INV_X1 U249 ( .A(n300), .ZN(n35) );
  OR2_X1 U250 ( .A1(n183), .A2(n151), .ZN(n285) );
  INV_X1 U251 ( .A(n87), .ZN(n286) );
  INV_X1 U252 ( .A(n319), .ZN(n287) );
  XOR2_X1 U253 ( .A(n245), .B(a[4]), .Z(n288) );
  XNOR2_X1 U254 ( .A(n115), .B(n305), .ZN(n289) );
  XNOR2_X1 U255 ( .A(n312), .B(b[7]), .ZN(n290) );
  CLKBUF_X3 U256 ( .A(n246), .Z(n312) );
  OR2_X1 U257 ( .A1(n46), .A2(n41), .ZN(n291) );
  CLKBUF_X1 U258 ( .A(n245), .Z(n292) );
  BUF_X2 U259 ( .A(n237), .Z(n334) );
  OAI21_X1 U260 ( .B1(n301), .B2(n47), .A(n42), .ZN(n293) );
  INV_X1 U261 ( .A(n243), .ZN(n294) );
  CLKBUF_X1 U262 ( .A(n25), .Z(n295) );
  XNOR2_X1 U263 ( .A(n247), .B(a[2]), .ZN(n296) );
  OAI22_X1 U264 ( .A1(n337), .A2(n203), .B1(n202), .B2(n333), .ZN(n297) );
  OAI22_X1 U265 ( .A1(n337), .A2(n203), .B1(n290), .B2(n333), .ZN(n110) );
  NOR2_X1 U266 ( .A1(n25), .A2(n20), .ZN(n298) );
  CLKBUF_X1 U267 ( .A(n59), .Z(n299) );
  NOR2_X1 U268 ( .A1(n125), .A2(n128), .ZN(n59) );
  CLKBUF_X1 U269 ( .A(n296), .Z(n323) );
  AND2_X1 U270 ( .A1(n102), .A2(n99), .ZN(n300) );
  NOR2_X1 U271 ( .A1(n103), .A2(n106), .ZN(n301) );
  AOI21_X1 U272 ( .B1(n331), .B2(n66), .A(n63), .ZN(n302) );
  OAI21_X2 U273 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  CLKBUF_X1 U274 ( .A(n47), .Z(n303) );
  CLKBUF_X1 U275 ( .A(n245), .Z(n304) );
  XNOR2_X1 U276 ( .A(n115), .B(n305), .ZN(n113) );
  XNOR2_X1 U277 ( .A(n120), .B(n117), .ZN(n305) );
  CLKBUF_X1 U278 ( .A(n300), .Z(n306) );
  INV_X1 U279 ( .A(n247), .ZN(n307) );
  INV_X2 U280 ( .A(n307), .ZN(n308) );
  NAND2_X1 U281 ( .A1(n115), .A2(n120), .ZN(n309) );
  NAND2_X1 U282 ( .A1(n115), .A2(n117), .ZN(n310) );
  NAND2_X1 U283 ( .A1(n120), .A2(n117), .ZN(n311) );
  NAND3_X1 U284 ( .A1(n309), .A2(n310), .A3(n311), .ZN(n112) );
  BUF_X1 U285 ( .A(n238), .Z(n333) );
  CLKBUF_X1 U286 ( .A(n56), .Z(n313) );
  CLKBUF_X1 U287 ( .A(n338), .Z(n314) );
  XOR2_X1 U288 ( .A(n244), .B(a[6]), .Z(n315) );
  XNOR2_X1 U289 ( .A(n245), .B(a[6]), .ZN(n316) );
  NAND2_X2 U290 ( .A1(n231), .A2(n255), .ZN(n235) );
  AOI21_X1 U291 ( .B1(n58), .B2(n50), .A(n51), .ZN(n339) );
  CLKBUF_X3 U292 ( .A(n227), .Z(n344) );
  XNOR2_X1 U293 ( .A(n31), .B(n317), .ZN(product[12]) );
  AND2_X1 U294 ( .A1(n328), .A2(n30), .ZN(n317) );
  NOR2_X1 U295 ( .A1(n113), .A2(n118), .ZN(n318) );
  NAND2_X1 U296 ( .A1(n244), .A2(b[1]), .ZN(n321) );
  NAND2_X1 U297 ( .A1(n319), .A2(n320), .ZN(n322) );
  NAND2_X1 U298 ( .A1(n321), .A2(n322), .ZN(n190) );
  INV_X1 U299 ( .A(n244), .ZN(n319) );
  INV_X1 U300 ( .A(b[1]), .ZN(n320) );
  NAND2_X1 U301 ( .A1(n230), .A2(n296), .ZN(n324) );
  AOI21_X1 U302 ( .B1(n306), .B2(n328), .A(n28), .ZN(n325) );
  NAND2_X1 U303 ( .A1(n288), .A2(n237), .ZN(n326) );
  INV_X1 U304 ( .A(n336), .ZN(n327) );
  XNOR2_X1 U305 ( .A(n48), .B(n5), .ZN(product[9]) );
  INV_X1 U306 ( .A(n293), .ZN(n38) );
  INV_X1 U307 ( .A(n46), .ZN(n85) );
  INV_X1 U308 ( .A(n295), .ZN(n23) );
  INV_X1 U309 ( .A(n77), .ZN(n75) );
  NOR2_X1 U310 ( .A1(n107), .A2(n112), .ZN(n46) );
  NAND2_X1 U311 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U312 ( .A(n41), .ZN(n84) );
  NAND2_X1 U313 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U314 ( .A(n299), .ZN(n88) );
  AOI21_X1 U315 ( .B1(n300), .B2(n328), .A(n28), .ZN(n26) );
  INV_X1 U316 ( .A(n30), .ZN(n28) );
  NAND2_X1 U317 ( .A1(n331), .A2(n65), .ZN(n9) );
  XOR2_X1 U318 ( .A(n22), .B(n1), .Z(product[13]) );
  NAND2_X1 U319 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U320 ( .A(n20), .ZN(n81) );
  XOR2_X1 U321 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U322 ( .A1(n87), .A2(n313), .ZN(n7) );
  INV_X1 U323 ( .A(n55), .ZN(n87) );
  XNOR2_X1 U324 ( .A(n54), .B(n6), .ZN(product[8]) );
  OAI21_X1 U325 ( .B1(n57), .B2(n286), .A(n313), .ZN(n54) );
  XNOR2_X1 U326 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U327 ( .A1(n330), .A2(n77), .ZN(n12) );
  NOR2_X1 U328 ( .A1(n46), .A2(n41), .ZN(n39) );
  NAND2_X1 U329 ( .A1(n329), .A2(n328), .ZN(n25) );
  OR2_X1 U330 ( .A1(n98), .A2(n97), .ZN(n328) );
  NOR2_X1 U331 ( .A1(n103), .A2(n106), .ZN(n41) );
  NAND2_X1 U332 ( .A1(n119), .A2(n124), .ZN(n56) );
  NOR2_X1 U333 ( .A1(n119), .A2(n124), .ZN(n55) );
  NAND2_X1 U334 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U335 ( .A(n71), .ZN(n91) );
  INV_X1 U336 ( .A(n94), .ZN(n95) );
  OR2_X1 U337 ( .A1(n169), .A2(n157), .ZN(n116) );
  XNOR2_X1 U338 ( .A(n169), .B(n157), .ZN(n117) );
  NOR2_X1 U339 ( .A1(n96), .A2(n95), .ZN(n20) );
  XOR2_X1 U340 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U341 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U342 ( .A(n67), .ZN(n90) );
  OR2_X1 U343 ( .A1(n99), .A2(n102), .ZN(n329) );
  NAND2_X1 U344 ( .A1(n125), .A2(n128), .ZN(n60) );
  INV_X1 U345 ( .A(n80), .ZN(n78) );
  INV_X1 U346 ( .A(n70), .ZN(n69) );
  NAND2_X1 U347 ( .A1(n98), .A2(n97), .ZN(n30) );
  NAND2_X1 U348 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U349 ( .A1(n182), .A2(n175), .ZN(n330) );
  NAND2_X1 U350 ( .A1(n103), .A2(n106), .ZN(n42) );
  OR2_X1 U351 ( .A1(n129), .A2(n132), .ZN(n331) );
  AND2_X1 U352 ( .A1(n344), .A2(n143), .ZN(n175) );
  INV_X1 U353 ( .A(n14), .ZN(product[15]) );
  OAI22_X1 U354 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  AND2_X1 U355 ( .A1(n344), .A2(n140), .ZN(n167) );
  OAI22_X1 U356 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  AND2_X1 U357 ( .A1(n344), .A2(n336), .ZN(n159) );
  OAI22_X1 U358 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OR2_X1 U359 ( .A1(n344), .A2(n241), .ZN(n201) );
  INV_X1 U360 ( .A(n100), .ZN(n101) );
  NOR2_X1 U361 ( .A1(n133), .A2(n134), .ZN(n67) );
  OAI22_X1 U362 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  INV_X1 U363 ( .A(n110), .ZN(n111) );
  NAND2_X1 U364 ( .A1(n135), .A2(n150), .ZN(n72) );
  INV_X1 U365 ( .A(n136), .ZN(n152) );
  NAND2_X1 U366 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U367 ( .A1(n341), .A2(n342), .ZN(n158) );
  OR2_X1 U368 ( .A1(n344), .A2(n240), .ZN(n192) );
  AND2_X1 U369 ( .A1(n285), .A2(n80), .ZN(product[1]) );
  XNOR2_X1 U370 ( .A(n245), .B(a[6]), .ZN(n236) );
  OR2_X1 U371 ( .A1(n344), .A2(n242), .ZN(n210) );
  INV_X1 U372 ( .A(n146), .ZN(n255) );
  OAI22_X1 U373 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OR2_X1 U374 ( .A1(n344), .A2(n243), .ZN(n219) );
  NAND2_X1 U375 ( .A1(n229), .A2(n237), .ZN(n233) );
  AND2_X1 U376 ( .A1(n344), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U377 ( .A(n287), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U378 ( .A(n287), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U379 ( .A(n287), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U380 ( .A(n287), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U381 ( .A(n244), .B(b[3]), .ZN(n188) );
  INV_X1 U382 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U383 ( .A(n247), .B(a[2]), .ZN(n238) );
  NOR2_X1 U384 ( .A1(n135), .A2(n150), .ZN(n71) );
  XNOR2_X1 U385 ( .A(n246), .B(a[4]), .ZN(n237) );
  INV_X1 U386 ( .A(n145), .ZN(n176) );
  OAI22_X1 U387 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  NAND2_X1 U388 ( .A1(n315), .A2(n236), .ZN(n335) );
  XOR2_X1 U389 ( .A(n245), .B(a[6]), .Z(n336) );
  NAND2_X1 U390 ( .A1(n228), .A2(n236), .ZN(n232) );
  XOR2_X1 U391 ( .A(n244), .B(a[6]), .Z(n228) );
  NAND2_X1 U392 ( .A1(n329), .A2(n35), .ZN(n3) );
  XOR2_X1 U393 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U394 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  AOI21_X1 U395 ( .B1(n330), .B2(n78), .A(n75), .ZN(n73) );
  NAND2_X1 U396 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U397 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  NAND2_X1 U398 ( .A1(n230), .A2(n238), .ZN(n337) );
  NAND2_X1 U399 ( .A1(n230), .A2(n296), .ZN(n234) );
  NOR2_X1 U400 ( .A1(n25), .A2(n20), .ZN(n18) );
  OAI21_X1 U401 ( .B1(n339), .B2(n291), .A(n38), .ZN(n338) );
  OAI21_X1 U402 ( .B1(n339), .B2(n291), .A(n38), .ZN(n36) );
  NAND2_X1 U403 ( .A1(n340), .A2(n53), .ZN(n6) );
  AOI21_X1 U404 ( .B1(n50), .B2(n58), .A(n51), .ZN(n49) );
  OR2_X1 U405 ( .A1(n289), .A2(n118), .ZN(n340) );
  NOR2_X1 U406 ( .A1(n232), .A2(n191), .ZN(n341) );
  NOR2_X1 U407 ( .A1(n190), .A2(n316), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n344), .B(n244), .ZN(n191) );
  INV_X1 U409 ( .A(n303), .ZN(n45) );
  OAI21_X1 U410 ( .B1(n301), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U411 ( .A1(n85), .A2(n303), .ZN(n5) );
  NAND2_X1 U412 ( .A1(n107), .A2(n112), .ZN(n47) );
  OAI21_X1 U413 ( .B1(n299), .B2(n302), .A(n60), .ZN(n343) );
  OAI21_X1 U414 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  INV_X1 U415 ( .A(n139), .ZN(n160) );
  XNOR2_X1 U416 ( .A(n244), .B(b[2]), .ZN(n189) );
  AOI21_X1 U417 ( .B1(n331), .B2(n66), .A(n63), .ZN(n61) );
  XNOR2_X1 U418 ( .A(n9), .B(n66), .ZN(product[5]) );
  INV_X1 U419 ( .A(n325), .ZN(n24) );
  OAI21_X1 U420 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  INV_X1 U421 ( .A(n142), .ZN(n168) );
  INV_X1 U422 ( .A(n343), .ZN(n57) );
  NAND2_X1 U423 ( .A1(n129), .A2(n132), .ZN(n65) );
  OAI22_X1 U424 ( .A1(n326), .A2(n199), .B1(n198), .B2(n334), .ZN(n165) );
  OAI22_X1 U425 ( .A1(n326), .A2(n197), .B1(n196), .B2(n334), .ZN(n163) );
  OAI22_X1 U426 ( .A1(n326), .A2(n194), .B1(n193), .B2(n334), .ZN(n100) );
  OAI22_X1 U427 ( .A1(n193), .A2(n326), .B1(n193), .B2(n334), .ZN(n139) );
  INV_X1 U428 ( .A(n334), .ZN(n140) );
  OAI22_X1 U429 ( .A1(n326), .A2(n196), .B1(n195), .B2(n334), .ZN(n162) );
  OAI22_X1 U430 ( .A1(n326), .A2(n198), .B1(n197), .B2(n334), .ZN(n164) );
  OAI22_X1 U431 ( .A1(n233), .A2(n195), .B1(n194), .B2(n334), .ZN(n161) );
  OAI22_X1 U432 ( .A1(n233), .A2(n241), .B1(n201), .B2(n334), .ZN(n149) );
  OAI22_X1 U433 ( .A1(n233), .A2(n200), .B1(n199), .B2(n334), .ZN(n166) );
  NAND2_X1 U434 ( .A1(n39), .A2(n298), .ZN(n16) );
  AOI21_X1 U435 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U436 ( .A(n8), .B(n302), .Z(product[6]) );
  OAI22_X1 U437 ( .A1(n184), .A2(n335), .B1(n184), .B2(n327), .ZN(n136) );
  NOR2_X1 U438 ( .A1(n52), .A2(n55), .ZN(n50) );
  OAI21_X1 U439 ( .B1(n318), .B2(n56), .A(n53), .ZN(n51) );
  NAND2_X1 U440 ( .A1(n289), .A2(n118), .ZN(n53) );
  NOR2_X1 U441 ( .A1(n113), .A2(n118), .ZN(n52) );
  OAI22_X1 U442 ( .A1(n335), .A2(n185), .B1(n184), .B2(n327), .ZN(n94) );
  OAI22_X1 U443 ( .A1(n335), .A2(n188), .B1(n187), .B2(n327), .ZN(n155) );
  OAI22_X1 U444 ( .A1(n335), .A2(n187), .B1(n186), .B2(n327), .ZN(n154) );
  OAI22_X1 U445 ( .A1(n335), .A2(n186), .B1(n185), .B2(n327), .ZN(n153) );
  OAI22_X1 U446 ( .A1(n335), .A2(n190), .B1(n189), .B2(n327), .ZN(n157) );
  OAI22_X1 U447 ( .A1(n335), .A2(n189), .B1(n327), .B2(n188), .ZN(n156) );
  OAI22_X1 U448 ( .A1(n232), .A2(n240), .B1(n192), .B2(n316), .ZN(n148) );
  XNOR2_X1 U449 ( .A(n304), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U450 ( .A(n292), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U451 ( .A(n304), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U452 ( .A(n304), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U453 ( .A(n245), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U454 ( .A(n292), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U455 ( .A(n344), .B(n292), .ZN(n200) );
  INV_X1 U456 ( .A(n245), .ZN(n241) );
  XOR2_X1 U457 ( .A(n245), .B(a[4]), .Z(n229) );
  INV_X1 U458 ( .A(n65), .ZN(n63) );
  OAI22_X1 U459 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  XNOR2_X1 U460 ( .A(n312), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U461 ( .A(n312), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U462 ( .A(n312), .B(b[5]), .ZN(n204) );
  XNOR2_X1 U463 ( .A(n312), .B(b[2]), .ZN(n207) );
  INV_X1 U464 ( .A(n312), .ZN(n242) );
  XNOR2_X1 U465 ( .A(n312), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U466 ( .A(n312), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U467 ( .A(n344), .B(n312), .ZN(n209) );
  XOR2_X1 U468 ( .A(n246), .B(a[2]), .Z(n230) );
  XNOR2_X1 U469 ( .A(n245), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U470 ( .A(n312), .B(b[1]), .ZN(n208) );
  NAND2_X1 U471 ( .A1(n183), .A2(n151), .ZN(n80) );
  AOI21_X1 U472 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  XOR2_X1 U473 ( .A(n43), .B(n4), .Z(product[10]) );
  OAI22_X1 U474 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  XNOR2_X1 U475 ( .A(n314), .B(n3), .ZN(product[11]) );
  AOI21_X1 U476 ( .B1(n338), .B2(n329), .A(n306), .ZN(n31) );
  AOI21_X1 U477 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U478 ( .B1(n49), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U479 ( .A(n339), .ZN(n48) );
  OAI22_X1 U480 ( .A1(n234), .A2(n204), .B1(n203), .B2(n333), .ZN(n169) );
  OAI22_X1 U481 ( .A1(n324), .A2(n207), .B1(n206), .B2(n333), .ZN(n172) );
  OAI22_X1 U482 ( .A1(n324), .A2(n206), .B1(n205), .B2(n323), .ZN(n171) );
  OAI22_X1 U483 ( .A1(n234), .A2(n205), .B1(n204), .B2(n296), .ZN(n170) );
  OAI22_X1 U484 ( .A1(n324), .A2(n208), .B1(n207), .B2(n323), .ZN(n173) );
  OAI22_X1 U485 ( .A1(n324), .A2(n242), .B1(n210), .B2(n323), .ZN(n150) );
  XNOR2_X1 U486 ( .A(n308), .B(b[5]), .ZN(n213) );
  OAI22_X1 U487 ( .A1(n290), .A2(n337), .B1(n202), .B2(n333), .ZN(n142) );
  XNOR2_X1 U488 ( .A(n294), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U489 ( .A(n308), .B(b[4]), .ZN(n214) );
  INV_X1 U490 ( .A(n333), .ZN(n143) );
  OAI22_X1 U491 ( .A1(n234), .A2(n209), .B1(n208), .B2(n296), .ZN(n174) );
  XNOR2_X1 U492 ( .A(n294), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U493 ( .A(n344), .B(n308), .ZN(n218) );
  XNOR2_X1 U494 ( .A(n308), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U495 ( .A(n308), .B(b[2]), .ZN(n216) );
  INV_X1 U496 ( .A(n247), .ZN(n243) );
  XNOR2_X1 U497 ( .A(n308), .B(b[1]), .ZN(n217) );
  XOR2_X1 U498 ( .A(n247), .B(n146), .Z(n231) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n33, n35,
         n36, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86,
         n87, n88, n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n142, n143, n145, n146, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n240, n241, n242, n243, n244, n245, n246,
         n247, n255, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n340, n341, n342, n343, n344;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n168), .B(n161), .CI(n334), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n156), .B(n162), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n164), .B(n177), .CI(n170), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n171), .B(n159), .CI(n178), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n166), .B(n149), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n181), .B(n174), .CO(n134), .S(n135) );
  XNOR2_X1 U249 ( .A(n169), .B(n157), .ZN(n117) );
  OR2_X1 U250 ( .A1(n183), .A2(n151), .ZN(n285) );
  OR2_X1 U251 ( .A1(n46), .A2(n41), .ZN(n286) );
  CLKBUF_X1 U252 ( .A(n246), .Z(n287) );
  CLKBUF_X1 U253 ( .A(n246), .Z(n288) );
  NOR2_X1 U254 ( .A1(n103), .A2(n106), .ZN(n289) );
  NOR2_X1 U255 ( .A1(n103), .A2(n106), .ZN(n41) );
  AND2_X1 U256 ( .A1(n336), .A2(n290), .ZN(n18) );
  AND2_X1 U257 ( .A1(n337), .A2(n81), .ZN(n290) );
  NAND2_X1 U258 ( .A1(n316), .A2(n317), .ZN(n291) );
  CLKBUF_X1 U259 ( .A(n246), .Z(n292) );
  CLKBUF_X1 U260 ( .A(n329), .Z(n293) );
  INV_X1 U261 ( .A(n241), .ZN(n294) );
  NAND2_X1 U262 ( .A1(n231), .A2(n255), .ZN(n295) );
  NAND2_X1 U263 ( .A1(n231), .A2(n255), .ZN(n235) );
  AOI21_X1 U264 ( .B1(n338), .B2(n66), .A(n63), .ZN(n296) );
  XOR2_X1 U265 ( .A(n243), .B(b[6]), .Z(n212) );
  NOR2_X1 U266 ( .A1(n125), .A2(n128), .ZN(n297) );
  NOR2_X1 U267 ( .A1(n125), .A2(n128), .ZN(n59) );
  OAI21_X1 U268 ( .B1(n289), .B2(n47), .A(n42), .ZN(n298) );
  OAI21_X1 U269 ( .B1(n297), .B2(n296), .A(n60), .ZN(n299) );
  CLKBUF_X1 U270 ( .A(n55), .Z(n300) );
  CLKBUF_X1 U271 ( .A(n328), .Z(n301) );
  CLKBUF_X1 U272 ( .A(n246), .Z(n302) );
  CLKBUF_X1 U273 ( .A(n328), .Z(n303) );
  BUF_X2 U274 ( .A(n238), .Z(n340) );
  BUF_X2 U275 ( .A(n244), .Z(n304) );
  XNOR2_X1 U276 ( .A(n115), .B(n309), .ZN(n305) );
  CLKBUF_X1 U277 ( .A(n247), .Z(n306) );
  CLKBUF_X1 U278 ( .A(n296), .Z(n307) );
  CLKBUF_X1 U279 ( .A(n299), .Z(n308) );
  XNOR2_X1 U280 ( .A(n115), .B(n309), .ZN(n113) );
  XNOR2_X1 U281 ( .A(n120), .B(n117), .ZN(n309) );
  OAI21_X1 U282 ( .B1(n52), .B2(n56), .A(n53), .ZN(n310) );
  CLKBUF_X1 U283 ( .A(n245), .Z(n311) );
  CLKBUF_X1 U284 ( .A(n66), .Z(n312) );
  CLKBUF_X1 U285 ( .A(n247), .Z(n313) );
  NAND2_X1 U286 ( .A1(n246), .A2(n315), .ZN(n316) );
  NAND2_X1 U287 ( .A1(n314), .A2(a[2]), .ZN(n317) );
  NAND2_X1 U288 ( .A1(n316), .A2(n317), .ZN(n230) );
  INV_X1 U289 ( .A(n246), .ZN(n314) );
  INV_X1 U290 ( .A(a[2]), .ZN(n315) );
  NOR2_X1 U291 ( .A1(n25), .A2(n20), .ZN(n318) );
  INV_X1 U292 ( .A(n33), .ZN(n319) );
  XNOR2_X1 U293 ( .A(n247), .B(a[2]), .ZN(n320) );
  OR2_X2 U294 ( .A1(n98), .A2(n97), .ZN(n337) );
  INV_X1 U295 ( .A(n35), .ZN(n321) );
  NAND2_X1 U296 ( .A1(n115), .A2(n120), .ZN(n322) );
  NAND2_X1 U297 ( .A1(n115), .A2(n117), .ZN(n323) );
  NAND2_X1 U298 ( .A1(n120), .A2(n117), .ZN(n324) );
  NAND3_X1 U299 ( .A1(n322), .A2(n323), .A3(n324), .ZN(n112) );
  CLKBUF_X1 U300 ( .A(n245), .Z(n325) );
  BUF_X2 U301 ( .A(n227), .Z(n344) );
  OAI21_X2 U302 ( .B1(n49), .B2(n286), .A(n38), .ZN(n36) );
  XNOR2_X1 U303 ( .A(n245), .B(a[6]), .ZN(n326) );
  CLKBUF_X3 U304 ( .A(n236), .Z(n343) );
  AOI21_X1 U305 ( .B1(n58), .B2(n50), .A(n51), .ZN(n327) );
  NAND2_X1 U306 ( .A1(n237), .A2(n229), .ZN(n328) );
  NAND2_X1 U307 ( .A1(n291), .A2(n320), .ZN(n329) );
  NAND2_X1 U308 ( .A1(n291), .A2(n320), .ZN(n330) );
  NAND2_X1 U309 ( .A1(n230), .A2(n320), .ZN(n234) );
  NOR2_X1 U310 ( .A1(n305), .A2(n118), .ZN(n331) );
  CLKBUF_X1 U311 ( .A(n232), .Z(n332) );
  AOI21_X1 U312 ( .B1(n33), .B2(n337), .A(n28), .ZN(n333) );
  OAI22_X1 U313 ( .A1(n329), .A2(n203), .B1(n340), .B2(n202), .ZN(n334) );
  INV_X1 U314 ( .A(n298), .ZN(n38) );
  INV_X1 U315 ( .A(n46), .ZN(n85) );
  INV_X1 U316 ( .A(n30), .ZN(n28) );
  NOR2_X1 U317 ( .A1(n107), .A2(n112), .ZN(n46) );
  AOI21_X1 U318 ( .B1(n50), .B2(n299), .A(n310), .ZN(n49) );
  NOR2_X1 U319 ( .A1(n113), .A2(n118), .ZN(n52) );
  NAND2_X1 U320 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U321 ( .A(n71), .ZN(n91) );
  NAND2_X1 U322 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U323 ( .A(n297), .ZN(n88) );
  NAND2_X1 U324 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U325 ( .A(n20), .ZN(n81) );
  NAND2_X1 U326 ( .A1(n337), .A2(n30), .ZN(n2) );
  XOR2_X1 U327 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U328 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U329 ( .A(n67), .ZN(n90) );
  XOR2_X1 U330 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U331 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U332 ( .A(n300), .ZN(n87) );
  XOR2_X1 U333 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U334 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U335 ( .A(n289), .ZN(n84) );
  XNOR2_X1 U336 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U337 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U338 ( .B1(n57), .B2(n300), .A(n56), .ZN(n54) );
  NOR2_X1 U339 ( .A1(n46), .A2(n41), .ZN(n39) );
  XNOR2_X1 U340 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U341 ( .A1(n335), .A2(n77), .ZN(n12) );
  INV_X1 U342 ( .A(n35), .ZN(n33) );
  NOR2_X1 U343 ( .A1(n119), .A2(n124), .ZN(n55) );
  OR2_X1 U344 ( .A1(n182), .A2(n175), .ZN(n335) );
  INV_X1 U345 ( .A(n94), .ZN(n95) );
  NOR2_X1 U346 ( .A1(n96), .A2(n95), .ZN(n20) );
  NAND2_X1 U347 ( .A1(n119), .A2(n124), .ZN(n56) );
  OR2_X1 U348 ( .A1(n99), .A2(n102), .ZN(n336) );
  NOR2_X1 U349 ( .A1(n133), .A2(n134), .ZN(n67) );
  INV_X1 U350 ( .A(n80), .ZN(n78) );
  NAND2_X1 U351 ( .A1(n133), .A2(n134), .ZN(n68) );
  NAND2_X1 U352 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U353 ( .A1(n129), .A2(n132), .ZN(n338) );
  INV_X1 U354 ( .A(n14), .ZN(product[15]) );
  OR2_X1 U355 ( .A1(n344), .A2(n242), .ZN(n210) );
  AND2_X1 U356 ( .A1(n344), .A2(n140), .ZN(n167) );
  OR2_X1 U357 ( .A1(n344), .A2(n241), .ZN(n201) );
  INV_X1 U358 ( .A(n139), .ZN(n160) );
  AND2_X1 U359 ( .A1(n344), .A2(n137), .ZN(n159) );
  INV_X1 U360 ( .A(n100), .ZN(n101) );
  INV_X1 U361 ( .A(n136), .ZN(n152) );
  OR2_X1 U362 ( .A1(n344), .A2(n240), .ZN(n192) );
  AND2_X1 U363 ( .A1(n285), .A2(n80), .ZN(product[1]) );
  NAND2_X1 U364 ( .A1(n229), .A2(n237), .ZN(n233) );
  INV_X1 U365 ( .A(n146), .ZN(n255) );
  NAND2_X1 U366 ( .A1(n228), .A2(n326), .ZN(n232) );
  AND2_X1 U367 ( .A1(n344), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U368 ( .A(n247), .B(a[2]), .ZN(n238) );
  XNOR2_X1 U369 ( .A(n304), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U370 ( .A(n304), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U371 ( .A(n304), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U372 ( .A(n344), .B(n304), .ZN(n191) );
  INV_X1 U373 ( .A(n244), .ZN(n240) );
  XOR2_X1 U374 ( .A(n244), .B(a[6]), .Z(n228) );
  NAND2_X1 U375 ( .A1(n125), .A2(n128), .ZN(n60) );
  OR2_X1 U376 ( .A1(n344), .A2(n243), .ZN(n219) );
  INV_X1 U377 ( .A(n145), .ZN(n176) );
  OR2_X1 U378 ( .A1(n169), .A2(n157), .ZN(n116) );
  AND2_X1 U379 ( .A1(n344), .A2(n143), .ZN(n175) );
  XNOR2_X1 U380 ( .A(n246), .B(a[4]), .ZN(n341) );
  XNOR2_X1 U381 ( .A(n246), .B(a[4]), .ZN(n342) );
  XNOR2_X1 U382 ( .A(n246), .B(a[4]), .ZN(n237) );
  INV_X1 U383 ( .A(n25), .ZN(n23) );
  OAI21_X1 U384 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  AOI21_X1 U385 ( .B1(n338), .B2(n66), .A(n63), .ZN(n61) );
  NAND2_X1 U386 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U387 ( .A1(n295), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U388 ( .A1(n295), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OAI22_X1 U389 ( .A1(n295), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U390 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  OAI22_X1 U391 ( .A1(n295), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U392 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OAI22_X1 U393 ( .A1(n295), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U394 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  NAND2_X1 U395 ( .A1(n338), .A2(n65), .ZN(n9) );
  INV_X1 U396 ( .A(n65), .ZN(n63) );
  OAI21_X1 U397 ( .B1(n41), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U398 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U399 ( .A(n47), .ZN(n45) );
  XNOR2_X1 U400 ( .A(n245), .B(a[6]), .ZN(n236) );
  NAND2_X1 U401 ( .A1(n103), .A2(n106), .ZN(n42) );
  NAND2_X1 U402 ( .A1(n336), .A2(n319), .ZN(n3) );
  NAND2_X1 U403 ( .A1(n336), .A2(n337), .ZN(n25) );
  INV_X1 U404 ( .A(n110), .ZN(n111) );
  NAND2_X1 U405 ( .A1(n107), .A2(n112), .ZN(n47) );
  INV_X1 U406 ( .A(n142), .ZN(n168) );
  XNOR2_X1 U407 ( .A(n9), .B(n312), .ZN(product[5]) );
  OAI21_X1 U408 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  OAI21_X1 U409 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  XOR2_X1 U410 ( .A(n11), .B(n73), .Z(product[3]) );
  INV_X1 U411 ( .A(n70), .ZN(n69) );
  AOI21_X1 U412 ( .B1(n335), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U413 ( .A(n77), .ZN(n75) );
  OAI22_X1 U414 ( .A1(n295), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  NAND2_X1 U415 ( .A1(n98), .A2(n97), .ZN(n30) );
  NAND2_X1 U416 ( .A1(n129), .A2(n132), .ZN(n65) );
  OAI22_X1 U417 ( .A1(n303), .A2(n199), .B1(n198), .B2(n342), .ZN(n165) );
  OAI22_X1 U418 ( .A1(n301), .A2(n197), .B1(n196), .B2(n342), .ZN(n163) );
  OAI22_X1 U419 ( .A1(n301), .A2(n194), .B1(n193), .B2(n341), .ZN(n100) );
  OAI22_X1 U420 ( .A1(n328), .A2(n198), .B1(n197), .B2(n341), .ZN(n164) );
  OAI22_X1 U421 ( .A1(n328), .A2(n196), .B1(n195), .B2(n341), .ZN(n162) );
  OAI22_X1 U422 ( .A1(n328), .A2(n195), .B1(n194), .B2(n342), .ZN(n161) );
  INV_X1 U423 ( .A(n342), .ZN(n140) );
  OAI22_X1 U424 ( .A1(n193), .A2(n303), .B1(n193), .B2(n341), .ZN(n139) );
  INV_X1 U425 ( .A(n288), .ZN(n242) );
  XNOR2_X1 U426 ( .A(n292), .B(b[4]), .ZN(n205) );
  OAI22_X1 U427 ( .A1(n233), .A2(n241), .B1(n201), .B2(n341), .ZN(n149) );
  XNOR2_X1 U428 ( .A(n287), .B(b[5]), .ZN(n204) );
  OAI22_X1 U429 ( .A1(n233), .A2(n200), .B1(n199), .B2(n342), .ZN(n166) );
  XNOR2_X1 U430 ( .A(n302), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U431 ( .A(n344), .B(n292), .ZN(n209) );
  INV_X1 U432 ( .A(n331), .ZN(n86) );
  NOR2_X1 U433 ( .A1(n331), .A2(n55), .ZN(n50) );
  OAI22_X1 U434 ( .A1(n184), .A2(n332), .B1(n184), .B2(n343), .ZN(n136) );
  OAI21_X1 U435 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  OAI22_X1 U436 ( .A1(n332), .A2(n185), .B1(n184), .B2(n343), .ZN(n94) );
  OAI22_X1 U437 ( .A1(n332), .A2(n188), .B1(n187), .B2(n343), .ZN(n155) );
  OAI22_X1 U438 ( .A1(n232), .A2(n187), .B1(n186), .B2(n343), .ZN(n154) );
  OAI22_X1 U439 ( .A1(n232), .A2(n186), .B1(n185), .B2(n343), .ZN(n153) );
  OAI22_X1 U440 ( .A1(n232), .A2(n190), .B1(n189), .B2(n343), .ZN(n157) );
  INV_X1 U441 ( .A(n343), .ZN(n137) );
  OAI22_X1 U442 ( .A1(n232), .A2(n189), .B1(n188), .B2(n343), .ZN(n156) );
  OAI22_X1 U443 ( .A1(n232), .A2(n240), .B1(n192), .B2(n343), .ZN(n148) );
  OAI22_X1 U444 ( .A1(n232), .A2(n191), .B1(n190), .B2(n343), .ZN(n158) );
  XNOR2_X1 U445 ( .A(n325), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U446 ( .A(n311), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U447 ( .A(n311), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U448 ( .A(n344), .B(n311), .ZN(n200) );
  INV_X1 U449 ( .A(n245), .ZN(n241) );
  XOR2_X1 U450 ( .A(n245), .B(a[4]), .Z(n229) );
  INV_X1 U451 ( .A(n333), .ZN(n24) );
  OAI21_X1 U452 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  AOI21_X1 U453 ( .B1(n321), .B2(n337), .A(n28), .ZN(n26) );
  NAND2_X1 U454 ( .A1(n102), .A2(n99), .ZN(n35) );
  NAND2_X1 U455 ( .A1(n305), .A2(n118), .ZN(n53) );
  XOR2_X1 U456 ( .A(n22), .B(n1), .Z(product[13]) );
  INV_X1 U457 ( .A(n308), .ZN(n57) );
  NOR2_X1 U458 ( .A1(n135), .A2(n150), .ZN(n71) );
  NAND2_X1 U459 ( .A1(n135), .A2(n150), .ZN(n72) );
  XNOR2_X1 U460 ( .A(n313), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U461 ( .A(n313), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U462 ( .A(n344), .B(n306), .ZN(n218) );
  INV_X1 U463 ( .A(n247), .ZN(n243) );
  XOR2_X1 U464 ( .A(n247), .B(n146), .Z(n231) );
  XOR2_X1 U465 ( .A(n31), .B(n2), .Z(product[12]) );
  XNOR2_X1 U466 ( .A(n304), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U467 ( .A(n325), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U468 ( .A(n246), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U469 ( .A(n247), .B(b[7]), .ZN(n211) );
  NAND2_X1 U470 ( .A1(n39), .A2(n318), .ZN(n16) );
  AOI21_X1 U471 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XNOR2_X1 U472 ( .A(n288), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U473 ( .A(n304), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U474 ( .A(n311), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U475 ( .A(n306), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U476 ( .A(n287), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U477 ( .A(n325), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U478 ( .A(n304), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U479 ( .A(n306), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U480 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U481 ( .A(n8), .B(n307), .Z(product[6]) );
  AOI21_X1 U482 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  NAND2_X1 U483 ( .A1(n183), .A2(n151), .ZN(n80) );
  XNOR2_X1 U484 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U485 ( .A(n294), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U486 ( .A(n302), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U487 ( .A(n313), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U488 ( .A(n36), .B(n3), .ZN(product[11]) );
  AOI21_X1 U489 ( .B1(n36), .B2(n336), .A(n33), .ZN(n31) );
  AOI21_X1 U490 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U491 ( .B1(n327), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U492 ( .A(n327), .ZN(n48) );
  OAI22_X1 U493 ( .A1(n330), .A2(n204), .B1(n203), .B2(n340), .ZN(n169) );
  OAI22_X1 U494 ( .A1(n293), .A2(n207), .B1(n206), .B2(n340), .ZN(n172) );
  OAI22_X1 U495 ( .A1(n330), .A2(n206), .B1(n205), .B2(n340), .ZN(n171) );
  OAI22_X1 U496 ( .A1(n329), .A2(n205), .B1(n204), .B2(n340), .ZN(n170) );
  OAI22_X1 U497 ( .A1(n330), .A2(n208), .B1(n207), .B2(n340), .ZN(n173) );
  OAI22_X1 U498 ( .A1(n293), .A2(n242), .B1(n210), .B2(n340), .ZN(n150) );
  OAI22_X1 U499 ( .A1(n329), .A2(n203), .B1(n340), .B2(n202), .ZN(n110) );
  OAI22_X1 U500 ( .A1(n234), .A2(n202), .B1(n202), .B2(n238), .ZN(n142) );
  INV_X1 U501 ( .A(n340), .ZN(n143) );
  OAI22_X1 U502 ( .A1(n330), .A2(n209), .B1(n208), .B2(n340), .ZN(n174) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_10_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  AND2_X1 U106 ( .A1(n155), .A2(n71), .ZN(SUM[0]) );
  CLKBUF_X1 U107 ( .A(n51), .Z(n143) );
  AOI21_X1 U108 ( .B1(n143), .B2(n154), .A(n48), .ZN(n144) );
  AOI21_X1 U109 ( .B1(n35), .B2(n151), .A(n32), .ZN(n145) );
  CLKBUF_X1 U110 ( .A(n43), .Z(n146) );
  XNOR2_X1 U111 ( .A(n16), .B(n147), .ZN(SUM[15]) );
  XOR2_X1 U112 ( .A(B[15]), .B(A[15]), .Z(n147) );
  INV_X1 U113 ( .A(n34), .ZN(n32) );
  INV_X1 U114 ( .A(n58), .ZN(n56) );
  AOI21_X1 U115 ( .B1(n67), .B2(n149), .A(n64), .ZN(n62) );
  INV_X1 U116 ( .A(n66), .ZN(n64) );
  NAND2_X1 U117 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U118 ( .A(n36), .ZN(n78) );
  AOI21_X1 U119 ( .B1(n51), .B2(n154), .A(n48), .ZN(n46) );
  INV_X1 U120 ( .A(n50), .ZN(n48) );
  NAND2_X1 U121 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U122 ( .A(n28), .ZN(n76) );
  NAND2_X1 U123 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U124 ( .A(n52), .ZN(n82) );
  NAND2_X1 U125 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U126 ( .A(n44), .ZN(n80) );
  NAND2_X1 U127 ( .A1(n152), .A2(n26), .ZN(n3) );
  NAND2_X1 U128 ( .A1(n153), .A2(n20), .ZN(n2) );
  NAND2_X1 U129 ( .A1(n148), .A2(n42), .ZN(n7) );
  NAND2_X1 U130 ( .A1(n149), .A2(n66), .ZN(n13) );
  NAND2_X1 U131 ( .A1(n150), .A2(n58), .ZN(n11) );
  NAND2_X1 U132 ( .A1(n151), .A2(n34), .ZN(n5) );
  XOR2_X1 U133 ( .A(n62), .B(n12), .Z(SUM[3]) );
  NAND2_X1 U134 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U135 ( .A(n60), .ZN(n84) );
  NAND2_X1 U136 ( .A1(n86), .A2(n69), .ZN(n14) );
  XNOR2_X1 U137 ( .A(n143), .B(n9), .ZN(SUM[6]) );
  NAND2_X1 U138 ( .A1(n154), .A2(n50), .ZN(n9) );
  INV_X1 U139 ( .A(n42), .ZN(n40) );
  INV_X1 U140 ( .A(n20), .ZN(n18) );
  INV_X1 U141 ( .A(n26), .ZN(n24) );
  OR2_X1 U142 ( .A1(A[8]), .A2(B[8]), .ZN(n148) );
  OR2_X1 U143 ( .A1(A[2]), .A2(B[2]), .ZN(n149) );
  NOR2_X1 U144 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  NOR2_X1 U145 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U146 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U147 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NOR2_X1 U148 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NAND2_X1 U149 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U150 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U151 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U152 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U153 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U154 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  OR2_X1 U155 ( .A1(A[4]), .A2(B[4]), .ZN(n150) );
  OR2_X1 U156 ( .A1(A[10]), .A2(B[10]), .ZN(n151) );
  OR2_X1 U157 ( .A1(A[12]), .A2(B[12]), .ZN(n152) );
  OR2_X1 U158 ( .A1(A[14]), .A2(B[14]), .ZN(n153) );
  OR2_X1 U159 ( .A1(A[6]), .A2(B[6]), .ZN(n154) );
  NAND2_X1 U160 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U161 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U162 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  NAND2_X1 U163 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U164 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  OR2_X1 U165 ( .A1(A[0]), .A2(B[0]), .ZN(n155) );
  OAI21_X1 U166 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  XOR2_X1 U167 ( .A(n54), .B(n10), .Z(SUM[5]) );
  AOI21_X1 U168 ( .B1(n59), .B2(n150), .A(n56), .ZN(n54) );
  XNOR2_X1 U169 ( .A(n27), .B(n3), .ZN(SUM[12]) );
  AOI21_X1 U170 ( .B1(n146), .B2(n148), .A(n40), .ZN(n156) );
  XOR2_X1 U171 ( .A(n14), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U172 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  OAI21_X1 U173 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U174 ( .A(n146), .B(n7), .ZN(SUM[8]) );
  INV_X1 U175 ( .A(n68), .ZN(n86) );
  AOI21_X1 U176 ( .B1(n43), .B2(n148), .A(n40), .ZN(n38) );
  NOR2_X1 U177 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  XNOR2_X1 U178 ( .A(n67), .B(n13), .ZN(SUM[2]) );
  XOR2_X1 U179 ( .A(n156), .B(n6), .Z(SUM[9]) );
  XOR2_X1 U180 ( .A(n144), .B(n8), .Z(SUM[7]) );
  XOR2_X1 U181 ( .A(n145), .B(n4), .Z(SUM[11]) );
  AOI21_X1 U182 ( .B1(n35), .B2(n151), .A(n32), .ZN(n30) );
  XNOR2_X1 U183 ( .A(n35), .B(n5), .ZN(SUM[10]) );
  NAND2_X1 U184 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  OAI21_X1 U185 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  OAI21_X1 U186 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U187 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  OAI21_X1 U188 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  XNOR2_X1 U189 ( .A(n59), .B(n11), .ZN(SUM[4]) );
  XNOR2_X1 U190 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  AOI21_X1 U191 ( .B1(n21), .B2(n153), .A(n18), .ZN(n16) );
  INV_X1 U192 ( .A(n22), .ZN(n73) );
  NAND2_X1 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  AOI21_X1 U194 ( .B1(n27), .B2(n152), .A(n24), .ZN(n22) );
endmodule


module add_layer_WIDTH16_10 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_10_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_9_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n157, n158;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  OR2_X1 U106 ( .A1(A[0]), .A2(B[0]), .ZN(n142) );
  CLKBUF_X1 U107 ( .A(n51), .Z(n143) );
  CLKBUF_X1 U108 ( .A(n27), .Z(n144) );
  CLKBUF_X1 U109 ( .A(n35), .Z(n145) );
  AOI21_X1 U110 ( .B1(n35), .B2(n152), .A(n32), .ZN(n146) );
  AOI21_X1 U111 ( .B1(n143), .B2(n155), .A(n48), .ZN(n147) );
  XNOR2_X1 U112 ( .A(n16), .B(n148), .ZN(SUM[15]) );
  XOR2_X1 U113 ( .A(B[15]), .B(A[15]), .Z(n148) );
  INV_X1 U114 ( .A(n34), .ZN(n32) );
  INV_X1 U115 ( .A(n58), .ZN(n56) );
  OAI21_X1 U116 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  INV_X1 U117 ( .A(n42), .ZN(n40) );
  AOI21_X1 U118 ( .B1(n67), .B2(n149), .A(n64), .ZN(n62) );
  INV_X1 U119 ( .A(n66), .ZN(n64) );
  AOI21_X1 U120 ( .B1(n51), .B2(n155), .A(n48), .ZN(n46) );
  INV_X1 U121 ( .A(n50), .ZN(n48) );
  NAND2_X1 U122 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U123 ( .A(n36), .ZN(n78) );
  NAND2_X1 U124 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U125 ( .A(n28), .ZN(n76) );
  NAND2_X1 U126 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U127 ( .A(n60), .ZN(n84) );
  NAND2_X1 U128 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U129 ( .A(n52), .ZN(n82) );
  NAND2_X1 U130 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U131 ( .A(n44), .ZN(n80) );
  NAND2_X1 U132 ( .A1(n155), .A2(n50), .ZN(n9) );
  NAND2_X1 U133 ( .A1(n153), .A2(n26), .ZN(n3) );
  NAND2_X1 U134 ( .A1(n152), .A2(n34), .ZN(n5) );
  NAND2_X1 U135 ( .A1(n150), .A2(n42), .ZN(n7) );
  XOR2_X1 U136 ( .A(n14), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U137 ( .A1(n86), .A2(n69), .ZN(n14) );
  XNOR2_X1 U138 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  NAND2_X1 U139 ( .A1(n154), .A2(n20), .ZN(n2) );
  XNOR2_X1 U140 ( .A(n67), .B(n13), .ZN(SUM[2]) );
  NAND2_X1 U141 ( .A1(n149), .A2(n66), .ZN(n13) );
  NAND2_X1 U142 ( .A1(n151), .A2(n58), .ZN(n11) );
  INV_X1 U143 ( .A(n20), .ZN(n18) );
  NAND2_X1 U144 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  INV_X1 U145 ( .A(n26), .ZN(n24) );
  OR2_X1 U146 ( .A1(A[2]), .A2(B[2]), .ZN(n149) );
  NOR2_X1 U147 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  NOR2_X1 U148 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U150 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NOR2_X1 U151 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NAND2_X1 U152 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U153 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U154 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  NAND2_X1 U155 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U156 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U157 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U158 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  OR2_X1 U159 ( .A1(A[8]), .A2(B[8]), .ZN(n150) );
  OR2_X1 U160 ( .A1(A[4]), .A2(B[4]), .ZN(n151) );
  OR2_X1 U161 ( .A1(A[10]), .A2(B[10]), .ZN(n152) );
  OR2_X1 U162 ( .A1(A[12]), .A2(B[12]), .ZN(n153) );
  OR2_X1 U163 ( .A1(A[14]), .A2(B[14]), .ZN(n154) );
  OR2_X1 U164 ( .A1(A[6]), .A2(B[6]), .ZN(n155) );
  NAND2_X1 U165 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U166 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U167 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  NAND2_X1 U168 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U169 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  AND2_X1 U170 ( .A1(n142), .A2(n71), .ZN(SUM[0]) );
  INV_X1 U171 ( .A(n68), .ZN(n86) );
  NOR2_X1 U172 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  XOR2_X1 U173 ( .A(n54), .B(n10), .Z(SUM[5]) );
  OAI21_X1 U174 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  AOI21_X1 U175 ( .B1(n59), .B2(n151), .A(n56), .ZN(n54) );
  CLKBUF_X1 U176 ( .A(n38), .Z(n157) );
  CLKBUF_X1 U177 ( .A(n59), .Z(n158) );
  AOI21_X1 U178 ( .B1(n43), .B2(n150), .A(n40), .ZN(n38) );
  XNOR2_X1 U179 ( .A(n43), .B(n7), .ZN(SUM[8]) );
  OAI21_X1 U180 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  OAI21_X1 U181 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U182 ( .A(n145), .B(n5), .ZN(SUM[10]) );
  XNOR2_X1 U183 ( .A(n143), .B(n9), .ZN(SUM[6]) );
  XOR2_X1 U184 ( .A(n157), .B(n6), .Z(SUM[9]) );
  XOR2_X1 U185 ( .A(n147), .B(n8), .Z(SUM[7]) );
  AOI21_X1 U186 ( .B1(n35), .B2(n152), .A(n32), .ZN(n30) );
  OAI21_X1 U187 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  XNOR2_X1 U188 ( .A(n158), .B(n11), .ZN(SUM[4]) );
  INV_X1 U189 ( .A(n22), .ZN(n73) );
  XNOR2_X1 U190 ( .A(n144), .B(n3), .ZN(SUM[12]) );
  XOR2_X1 U191 ( .A(n62), .B(n12), .Z(SUM[3]) );
  AOI21_X1 U192 ( .B1(n27), .B2(n153), .A(n24), .ZN(n22) );
  OAI21_X1 U193 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  NAND2_X1 U194 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  AOI21_X1 U195 ( .B1(n21), .B2(n154), .A(n18), .ZN(n16) );
  XOR2_X1 U196 ( .A(n146), .B(n4), .Z(SUM[11]) );
endmodule


module add_layer_WIDTH16_9 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_9_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37,
         n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70,
         n71, n73, n75, n77, n79, n81, n82, n83, n84, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n71), .CO(n16), .S(SUM[14]) );
  OR2_X1 U104 ( .A1(A[0]), .A2(B[0]), .ZN(n140) );
  CLKBUF_X1 U105 ( .A(n22), .Z(n141) );
  CLKBUF_X1 U106 ( .A(n25), .Z(n142) );
  CLKBUF_X1 U107 ( .A(n66), .Z(n143) );
  AOI21_X1 U108 ( .B1(n58), .B2(n143), .A(n59), .ZN(n144) );
  CLKBUF_X1 U109 ( .A(n41), .Z(n145) );
  CLKBUF_X1 U110 ( .A(n54), .Z(n146) );
  CLKBUF_X1 U111 ( .A(n38), .Z(n147) );
  AOI21_X1 U112 ( .B1(n54), .B2(n153), .A(n51), .ZN(n148) );
  AOI21_X1 U113 ( .B1(n38), .B2(n156), .A(n35), .ZN(n149) );
  NOR2_X1 U114 ( .A1(A[3]), .A2(B[3]), .ZN(n150) );
  INV_X1 U115 ( .A(n29), .ZN(n27) );
  INV_X1 U116 ( .A(n45), .ZN(n43) );
  INV_X1 U117 ( .A(n53), .ZN(n51) );
  AOI21_X1 U118 ( .B1(n58), .B2(n66), .A(n59), .ZN(n57) );
  AOI21_X1 U119 ( .B1(n147), .B2(n156), .A(n35), .ZN(n33) );
  INV_X1 U120 ( .A(n37), .ZN(n35) );
  OAI21_X1 U121 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  NAND2_X1 U122 ( .A1(n79), .A2(n48), .ZN(n9) );
  INV_X1 U123 ( .A(n47), .ZN(n79) );
  NAND2_X1 U124 ( .A1(n77), .A2(n40), .ZN(n7) );
  INV_X1 U125 ( .A(n39), .ZN(n77) );
  NAND2_X1 U126 ( .A1(n156), .A2(n37), .ZN(n6) );
  XOR2_X1 U127 ( .A(n14), .B(n70), .Z(SUM[1]) );
  NAND2_X1 U128 ( .A1(n84), .A2(n68), .ZN(n14) );
  INV_X1 U129 ( .A(n67), .ZN(n84) );
  XOR2_X1 U130 ( .A(n65), .B(n13), .Z(SUM[2]) );
  INV_X1 U131 ( .A(n63), .ZN(n83) );
  XOR2_X1 U132 ( .A(n33), .B(n5), .Z(SUM[10]) );
  NAND2_X1 U133 ( .A1(n75), .A2(n32), .ZN(n5) );
  INV_X1 U134 ( .A(n31), .ZN(n75) );
  XOR2_X1 U135 ( .A(n144), .B(n11), .Z(SUM[4]) );
  NAND2_X1 U136 ( .A1(n81), .A2(n56), .ZN(n11) );
  INV_X1 U137 ( .A(n55), .ZN(n81) );
  NAND2_X1 U138 ( .A1(n152), .A2(n45), .ZN(n8) );
  NAND2_X1 U139 ( .A1(n153), .A2(n53), .ZN(n10) );
  XNOR2_X1 U140 ( .A(n62), .B(n12), .ZN(SUM[3]) );
  NAND2_X1 U141 ( .A1(n82), .A2(n61), .ZN(n12) );
  NAND2_X1 U142 ( .A1(n155), .A2(n29), .ZN(n4) );
  NAND2_X1 U143 ( .A1(n154), .A2(n21), .ZN(n2) );
  NAND2_X1 U144 ( .A1(n73), .A2(n24), .ZN(n3) );
  INV_X1 U145 ( .A(n23), .ZN(n73) );
  NOR2_X1 U146 ( .A1(A[2]), .A2(B[2]), .ZN(n63) );
  XNOR2_X1 U147 ( .A(n16), .B(n151), .ZN(SUM[15]) );
  XNOR2_X1 U148 ( .A(B[15]), .B(A[15]), .ZN(n151) );
  NOR2_X1 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U150 ( .A1(A[1]), .A2(B[1]), .ZN(n67) );
  NAND2_X1 U151 ( .A1(A[0]), .A2(B[0]), .ZN(n70) );
  NOR2_X1 U152 ( .A1(A[4]), .A2(B[4]), .ZN(n55) );
  NOR2_X1 U153 ( .A1(A[8]), .A2(B[8]), .ZN(n39) );
  NOR2_X1 U154 ( .A1(A[6]), .A2(B[6]), .ZN(n47) );
  NOR2_X1 U155 ( .A1(A[10]), .A2(B[10]), .ZN(n31) );
  NOR2_X1 U156 ( .A1(A[12]), .A2(B[12]), .ZN(n23) );
  INV_X1 U157 ( .A(n21), .ZN(n19) );
  NAND2_X1 U158 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U159 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U160 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U161 ( .A1(A[13]), .A2(B[13]), .ZN(n21) );
  NAND2_X1 U162 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U163 ( .A1(A[4]), .A2(B[4]), .ZN(n56) );
  OR2_X1 U164 ( .A1(A[7]), .A2(B[7]), .ZN(n152) );
  OR2_X1 U165 ( .A1(A[5]), .A2(B[5]), .ZN(n153) );
  OR2_X1 U166 ( .A1(A[13]), .A2(B[13]), .ZN(n154) );
  OR2_X1 U167 ( .A1(A[11]), .A2(B[11]), .ZN(n155) );
  OR2_X1 U168 ( .A1(A[9]), .A2(B[9]), .ZN(n156) );
  NAND2_X1 U169 ( .A1(A[8]), .A2(B[8]), .ZN(n40) );
  NAND2_X1 U170 ( .A1(A[6]), .A2(B[6]), .ZN(n48) );
  NAND2_X1 U171 ( .A1(A[10]), .A2(B[10]), .ZN(n32) );
  NAND2_X1 U172 ( .A1(A[12]), .A2(B[12]), .ZN(n24) );
  AND2_X1 U173 ( .A1(n140), .A2(n70), .ZN(SUM[0]) );
  NAND2_X1 U174 ( .A1(n83), .A2(n64), .ZN(n13) );
  OAI21_X1 U175 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  XNOR2_X1 U176 ( .A(n30), .B(n4), .ZN(SUM[11]) );
  XNOR2_X1 U177 ( .A(n46), .B(n8), .ZN(SUM[7]) );
  AOI21_X1 U178 ( .B1(n46), .B2(n152), .A(n43), .ZN(n41) );
  XOR2_X1 U179 ( .A(n145), .B(n7), .Z(SUM[8]) );
  OAI21_X1 U180 ( .B1(n148), .B2(n47), .A(n48), .ZN(n46) );
  XOR2_X1 U181 ( .A(n49), .B(n9), .Z(SUM[6]) );
  AOI21_X1 U182 ( .B1(n146), .B2(n153), .A(n51), .ZN(n49) );
  XNOR2_X1 U183 ( .A(n147), .B(n6), .ZN(SUM[9]) );
  XNOR2_X1 U184 ( .A(n146), .B(n10), .ZN(SUM[5]) );
  INV_X1 U185 ( .A(n143), .ZN(n65) );
  NAND2_X1 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n64) );
  OAI21_X1 U187 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U188 ( .B1(n67), .B2(n70), .A(n68), .ZN(n66) );
  AOI21_X1 U189 ( .B1(n30), .B2(n155), .A(n27), .ZN(n25) );
  OAI21_X1 U190 ( .B1(n149), .B2(n31), .A(n32), .ZN(n30) );
  NAND2_X1 U191 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  INV_X1 U192 ( .A(n17), .ZN(n71) );
  OAI21_X1 U193 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
  AOI21_X1 U194 ( .B1(n22), .B2(n154), .A(n19), .ZN(n17) );
  XOR2_X1 U195 ( .A(n142), .B(n3), .Z(SUM[12]) );
  XNOR2_X1 U196 ( .A(n141), .B(n2), .ZN(SUM[13]) );
  NAND2_X1 U197 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  OAI21_X1 U198 ( .B1(n60), .B2(n64), .A(n61), .ZN(n59) );
  NOR2_X1 U199 ( .A1(n63), .A2(n150), .ZN(n58) );
  INV_X1 U200 ( .A(n150), .ZN(n82) );
endmodule


module add_layer_WIDTH16_3 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_3_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_3 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_3 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_3 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_10 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_9 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_3 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_3 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12 \genblk1[0].mult  ( .clk(clk), 
        .ia({\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11 \genblk1[1].mult  ( .clk(clk), 
        .ia({\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10 \genblk1[2].mult  ( .clk(clk), 
        .ia({\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9 \genblk1[3].mult  ( .clk(clk), .ia(
        {\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_3 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n33, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n85, n86,
         n87, n88, n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n142, n143, n145, n146, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n240, n241, n242, n243, n244, n245, n246,
         n247, n255, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n168), .B(n110), .CI(n161), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n156), .B(n162), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n170), .B(n177), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n181), .B(n174), .CO(n134), .S(n135) );
  NOR2_X1 U249 ( .A1(n103), .A2(n106), .ZN(n41) );
  OR2_X1 U250 ( .A1(n183), .A2(n151), .ZN(n285) );
  INV_X1 U251 ( .A(n299), .ZN(n286) );
  OAI21_X1 U252 ( .B1(n41), .B2(n47), .A(n42), .ZN(n287) );
  CLKBUF_X1 U253 ( .A(n61), .Z(n288) );
  XOR2_X1 U254 ( .A(n241), .B(b[4]), .Z(n196) );
  OAI21_X1 U255 ( .B1(n59), .B2(n61), .A(n60), .ZN(n289) );
  NOR2_X2 U256 ( .A1(n125), .A2(n128), .ZN(n59) );
  OR2_X1 U257 ( .A1(n103), .A2(n106), .ZN(n290) );
  XNOR2_X1 U258 ( .A(n338), .B(b[7]), .ZN(n291) );
  CLKBUF_X1 U259 ( .A(n245), .Z(n292) );
  XNOR2_X1 U260 ( .A(n293), .B(n122), .ZN(n115) );
  XNOR2_X1 U261 ( .A(n163), .B(n176), .ZN(n293) );
  XNOR2_X1 U262 ( .A(a[2]), .B(n247), .ZN(n294) );
  NAND2_X2 U263 ( .A1(n231), .A2(n255), .ZN(n235) );
  INV_X2 U264 ( .A(n146), .ZN(n255) );
  INV_X1 U265 ( .A(n240), .ZN(n295) );
  XNOR2_X1 U266 ( .A(n338), .B(b[7]), .ZN(n296) );
  INV_X1 U267 ( .A(n143), .ZN(n297) );
  CLKBUF_X1 U268 ( .A(n55), .Z(n298) );
  NAND2_X1 U269 ( .A1(n244), .A2(n300), .ZN(n301) );
  NAND2_X1 U270 ( .A1(n299), .A2(a[6]), .ZN(n302) );
  NAND2_X1 U271 ( .A1(n301), .A2(n302), .ZN(n318) );
  INV_X1 U272 ( .A(n244), .ZN(n299) );
  INV_X1 U273 ( .A(a[6]), .ZN(n300) );
  NAND2_X2 U274 ( .A1(n318), .A2(n236), .ZN(n328) );
  OAI21_X1 U275 ( .B1(n67), .B2(n69), .A(n68), .ZN(n303) );
  CLKBUF_X1 U276 ( .A(n33), .Z(n304) );
  BUF_X1 U277 ( .A(n238), .Z(n341) );
  CLKBUF_X1 U278 ( .A(n56), .Z(n305) );
  XNOR2_X1 U279 ( .A(n306), .B(n115), .ZN(n113) );
  XNOR2_X1 U280 ( .A(n120), .B(n117), .ZN(n306) );
  CLKBUF_X3 U281 ( .A(n247), .Z(n336) );
  XOR2_X1 U282 ( .A(n172), .B(n179), .Z(n307) );
  XOR2_X1 U283 ( .A(n307), .B(n131), .Z(n129) );
  NAND2_X1 U284 ( .A1(n131), .A2(n172), .ZN(n308) );
  NAND2_X1 U285 ( .A1(n131), .A2(n179), .ZN(n309) );
  NAND2_X1 U286 ( .A1(n172), .A2(n179), .ZN(n310) );
  NAND3_X1 U287 ( .A1(n308), .A2(n309), .A3(n310), .ZN(n128) );
  NAND2_X1 U288 ( .A1(n163), .A2(n176), .ZN(n311) );
  NAND2_X1 U289 ( .A1(n163), .A2(n122), .ZN(n312) );
  NAND2_X1 U290 ( .A1(n176), .A2(n122), .ZN(n313) );
  NAND3_X1 U291 ( .A1(n311), .A2(n312), .A3(n313), .ZN(n114) );
  NAND2_X1 U292 ( .A1(n120), .A2(n117), .ZN(n314) );
  NAND2_X1 U293 ( .A1(n120), .A2(n115), .ZN(n315) );
  NAND2_X1 U294 ( .A1(n117), .A2(n115), .ZN(n316) );
  NAND3_X1 U295 ( .A1(n314), .A2(n315), .A3(n316), .ZN(n112) );
  CLKBUF_X1 U296 ( .A(n343), .Z(n317) );
  BUF_X2 U297 ( .A(n227), .Z(n343) );
  CLKBUF_X1 U298 ( .A(n245), .Z(n319) );
  BUF_X2 U299 ( .A(n246), .Z(n339) );
  OAI21_X2 U300 ( .B1(n342), .B2(n37), .A(n38), .ZN(n36) );
  BUF_X2 U301 ( .A(n246), .Z(n338) );
  NAND2_X1 U302 ( .A1(n229), .A2(n237), .ZN(n320) );
  NAND2_X1 U303 ( .A1(n245), .A2(n322), .ZN(n323) );
  NAND2_X1 U304 ( .A1(n321), .A2(a[4]), .ZN(n324) );
  NAND2_X1 U305 ( .A1(n323), .A2(n324), .ZN(n229) );
  INV_X1 U306 ( .A(n245), .ZN(n321) );
  INV_X1 U307 ( .A(a[4]), .ZN(n322) );
  NAND2_X1 U308 ( .A1(n229), .A2(n237), .ZN(n233) );
  XNOR2_X2 U309 ( .A(n339), .B(a[4]), .ZN(n337) );
  AOI21_X1 U310 ( .B1(n304), .B2(n329), .A(n28), .ZN(n325) );
  INV_X1 U311 ( .A(n143), .ZN(n326) );
  NOR2_X1 U312 ( .A1(n113), .A2(n118), .ZN(n327) );
  XOR2_X1 U313 ( .A(n246), .B(a[2]), .Z(n230) );
  NAND2_X1 U314 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U315 ( .A(n46), .ZN(n85) );
  INV_X1 U316 ( .A(n25), .ZN(n23) );
  INV_X1 U317 ( .A(n47), .ZN(n45) );
  INV_X1 U318 ( .A(n287), .ZN(n38) );
  INV_X1 U319 ( .A(n39), .ZN(n37) );
  INV_X1 U320 ( .A(n77), .ZN(n75) );
  NOR2_X1 U321 ( .A1(n107), .A2(n112), .ZN(n46) );
  INV_X1 U322 ( .A(n70), .ZN(n69) );
  NAND2_X1 U323 ( .A1(n107), .A2(n112), .ZN(n47) );
  OAI21_X1 U324 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  OAI21_X1 U325 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  NOR2_X1 U326 ( .A1(n113), .A2(n118), .ZN(n52) );
  AOI21_X1 U327 ( .B1(n330), .B2(n66), .A(n63), .ZN(n61) );
  INV_X1 U328 ( .A(n65), .ZN(n63) );
  NAND2_X1 U329 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U330 ( .A(n20), .ZN(n81) );
  NAND2_X1 U331 ( .A1(n329), .A2(n30), .ZN(n2) );
  AOI21_X1 U332 ( .B1(n33), .B2(n329), .A(n28), .ZN(n26) );
  INV_X1 U333 ( .A(n30), .ZN(n28) );
  XOR2_X1 U334 ( .A(n11), .B(n73), .Z(product[3]) );
  INV_X1 U335 ( .A(n71), .ZN(n91) );
  XOR2_X1 U336 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U337 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U338 ( .A(n67), .ZN(n90) );
  XOR2_X1 U339 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U340 ( .A1(n290), .A2(n42), .ZN(n4) );
  XOR2_X1 U341 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U342 ( .A1(n87), .A2(n305), .ZN(n7) );
  INV_X1 U343 ( .A(n298), .ZN(n87) );
  OAI21_X1 U344 ( .B1(n41), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U345 ( .A1(n113), .A2(n118), .ZN(n53) );
  XNOR2_X1 U346 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U347 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U348 ( .B1(n57), .B2(n298), .A(n305), .ZN(n54) );
  XNOR2_X1 U349 ( .A(n9), .B(n303), .ZN(product[5]) );
  NAND2_X1 U350 ( .A1(n330), .A2(n65), .ZN(n9) );
  XNOR2_X1 U351 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U352 ( .A1(n331), .A2(n77), .ZN(n12) );
  NOR2_X1 U353 ( .A1(n46), .A2(n41), .ZN(n39) );
  NOR2_X1 U354 ( .A1(n25), .A2(n20), .ZN(n18) );
  INV_X1 U355 ( .A(n35), .ZN(n33) );
  NAND2_X1 U356 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U357 ( .A(n59), .ZN(n88) );
  OR2_X1 U358 ( .A1(n169), .A2(n157), .ZN(n116) );
  NOR2_X1 U359 ( .A1(n133), .A2(n134), .ZN(n67) );
  NOR2_X1 U360 ( .A1(n96), .A2(n95), .ZN(n20) );
  NOR2_X1 U361 ( .A1(n119), .A2(n124), .ZN(n55) );
  XNOR2_X1 U362 ( .A(n169), .B(n157), .ZN(n117) );
  OR2_X1 U363 ( .A1(n98), .A2(n97), .ZN(n329) );
  INV_X1 U364 ( .A(n94), .ZN(n95) );
  OR2_X1 U365 ( .A1(n129), .A2(n132), .ZN(n330) );
  NAND2_X1 U366 ( .A1(n119), .A2(n124), .ZN(n56) );
  NAND2_X1 U367 ( .A1(n103), .A2(n106), .ZN(n42) );
  NAND2_X1 U368 ( .A1(n125), .A2(n128), .ZN(n60) );
  INV_X1 U369 ( .A(n80), .ZN(n78) );
  NAND2_X1 U370 ( .A1(n98), .A2(n97), .ZN(n30) );
  NAND2_X1 U371 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U372 ( .A1(n182), .A2(n175), .ZN(n331) );
  OR2_X1 U373 ( .A1(n99), .A2(n102), .ZN(n332) );
  INV_X1 U374 ( .A(n14), .ZN(product[15]) );
  OR2_X1 U375 ( .A1(n343), .A2(n242), .ZN(n210) );
  OR2_X1 U376 ( .A1(n343), .A2(n241), .ZN(n201) );
  AND2_X1 U377 ( .A1(n343), .A2(n137), .ZN(n159) );
  OAI22_X1 U378 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  INV_X1 U379 ( .A(n100), .ZN(n101) );
  AND2_X1 U380 ( .A1(n317), .A2(n140), .ZN(n167) );
  OAI22_X1 U381 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  INV_X1 U382 ( .A(n142), .ZN(n168) );
  OAI22_X1 U383 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  INV_X1 U384 ( .A(n136), .ZN(n152) );
  OR2_X1 U385 ( .A1(n343), .A2(n240), .ZN(n192) );
  INV_X1 U386 ( .A(n145), .ZN(n176) );
  AND2_X1 U387 ( .A1(n285), .A2(n80), .ZN(product[1]) );
  AND2_X1 U388 ( .A1(n343), .A2(n143), .ZN(n175) );
  XNOR2_X1 U389 ( .A(n247), .B(a[2]), .ZN(n238) );
  OAI22_X1 U390 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OR2_X1 U391 ( .A1(n343), .A2(n243), .ZN(n219) );
  NAND2_X1 U392 ( .A1(n228), .A2(n335), .ZN(n232) );
  AND2_X1 U393 ( .A1(n317), .A2(n146), .ZN(product[0]) );
  NOR2_X1 U394 ( .A1(n135), .A2(n150), .ZN(n71) );
  NAND2_X1 U395 ( .A1(n133), .A2(n134), .ZN(n68) );
  XNOR2_X1 U396 ( .A(n245), .B(a[6]), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n245), .B(a[6]), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n245), .B(a[6]), .ZN(n236) );
  NAND2_X1 U399 ( .A1(n129), .A2(n132), .ZN(n65) );
  XNOR2_X1 U400 ( .A(n295), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U401 ( .A(n295), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U402 ( .A(n295), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U403 ( .A(n286), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U404 ( .A(n343), .B(n286), .ZN(n191) );
  INV_X1 U405 ( .A(n244), .ZN(n240) );
  XOR2_X1 U406 ( .A(n244), .B(a[6]), .Z(n228) );
  OAI22_X1 U407 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  NAND2_X1 U408 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U409 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  INV_X1 U410 ( .A(n325), .ZN(n24) );
  OAI21_X1 U411 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  INV_X1 U412 ( .A(n110), .ZN(n111) );
  XNOR2_X1 U413 ( .A(n295), .B(b[6]), .ZN(n185) );
  OAI22_X1 U414 ( .A1(n216), .A2(n235), .B1(n215), .B2(n255), .ZN(n181) );
  OAI22_X1 U415 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U416 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  XNOR2_X1 U417 ( .A(n339), .B(a[4]), .ZN(n237) );
  XNOR2_X1 U418 ( .A(n286), .B(b[2]), .ZN(n189) );
  NAND2_X1 U419 ( .A1(n230), .A2(n294), .ZN(n340) );
  NAND2_X1 U420 ( .A1(n230), .A2(n294), .ZN(n234) );
  NAND2_X1 U421 ( .A1(n183), .A2(n151), .ZN(n80) );
  INV_X1 U422 ( .A(n327), .ZN(n86) );
  NOR2_X1 U423 ( .A1(n327), .A2(n55), .ZN(n50) );
  OAI21_X1 U424 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  INV_X1 U425 ( .A(n139), .ZN(n160) );
  AOI21_X1 U426 ( .B1(n331), .B2(n78), .A(n75), .ZN(n73) );
  AOI21_X1 U427 ( .B1(n50), .B2(n289), .A(n51), .ZN(n342) );
  AOI21_X1 U428 ( .B1(n50), .B2(n58), .A(n51), .ZN(n49) );
  OAI21_X1 U429 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  NAND2_X1 U430 ( .A1(n91), .A2(n72), .ZN(n11) );
  NAND2_X1 U431 ( .A1(n332), .A2(n35), .ZN(n3) );
  NAND2_X1 U432 ( .A1(n332), .A2(n329), .ZN(n25) );
  NAND2_X1 U433 ( .A1(n102), .A2(n99), .ZN(n35) );
  XOR2_X1 U434 ( .A(n22), .B(n1), .Z(product[13]) );
  OAI22_X1 U435 ( .A1(n184), .A2(n328), .B1(n184), .B2(n334), .ZN(n136) );
  OAI22_X1 U436 ( .A1(n328), .A2(n185), .B1(n184), .B2(n335), .ZN(n94) );
  OAI22_X1 U437 ( .A1(n328), .A2(n188), .B1(n187), .B2(n334), .ZN(n155) );
  OAI22_X1 U438 ( .A1(n328), .A2(n187), .B1(n186), .B2(n334), .ZN(n154) );
  OAI22_X1 U439 ( .A1(n328), .A2(n186), .B1(n185), .B2(n334), .ZN(n153) );
  INV_X1 U440 ( .A(n334), .ZN(n137) );
  OAI22_X1 U441 ( .A1(n328), .A2(n190), .B1(n189), .B2(n335), .ZN(n157) );
  OAI22_X1 U442 ( .A1(n189), .A2(n328), .B1(n188), .B2(n335), .ZN(n156) );
  XNOR2_X1 U443 ( .A(n319), .B(b[2]), .ZN(n198) );
  OAI22_X1 U444 ( .A1(n232), .A2(n240), .B1(n192), .B2(n335), .ZN(n148) );
  OAI22_X1 U445 ( .A1(n232), .A2(n191), .B1(n190), .B2(n334), .ZN(n158) );
  XNOR2_X1 U446 ( .A(n319), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U447 ( .A(n319), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U448 ( .A(n343), .B(n292), .ZN(n200) );
  XNOR2_X1 U449 ( .A(n292), .B(b[5]), .ZN(n195) );
  INV_X1 U450 ( .A(n245), .ZN(n241) );
  XNOR2_X1 U451 ( .A(n245), .B(b[6]), .ZN(n194) );
  NAND2_X1 U452 ( .A1(n39), .A2(n18), .ZN(n16) );
  AOI21_X1 U453 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U454 ( .A(n31), .B(n2), .Z(product[12]) );
  INV_X1 U455 ( .A(n289), .ZN(n57) );
  NAND2_X1 U456 ( .A1(n135), .A2(n150), .ZN(n72) );
  XNOR2_X1 U457 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U458 ( .A(n8), .B(n288), .Z(product[6]) );
  AOI21_X1 U459 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  OAI22_X1 U460 ( .A1(n320), .A2(n199), .B1(n198), .B2(n337), .ZN(n165) );
  OAI22_X1 U461 ( .A1(n320), .A2(n197), .B1(n196), .B2(n337), .ZN(n163) );
  OAI22_X1 U462 ( .A1(n320), .A2(n194), .B1(n193), .B2(n337), .ZN(n100) );
  OAI22_X1 U463 ( .A1(n233), .A2(n196), .B1(n195), .B2(n337), .ZN(n162) );
  OAI22_X1 U464 ( .A1(n320), .A2(n198), .B1(n197), .B2(n337), .ZN(n164) );
  OAI22_X1 U465 ( .A1(n193), .A2(n320), .B1(n193), .B2(n337), .ZN(n139) );
  OAI22_X1 U466 ( .A1(n233), .A2(n195), .B1(n194), .B2(n337), .ZN(n161) );
  INV_X1 U467 ( .A(n337), .ZN(n140) );
  OAI22_X1 U468 ( .A1(n233), .A2(n241), .B1(n201), .B2(n337), .ZN(n149) );
  XNOR2_X1 U469 ( .A(n338), .B(b[3]), .ZN(n206) );
  OAI22_X1 U470 ( .A1(n233), .A2(n200), .B1(n199), .B2(n337), .ZN(n166) );
  XNOR2_X1 U471 ( .A(n338), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U472 ( .A(n338), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U473 ( .A(n338), .B(b[5]), .ZN(n204) );
  INV_X1 U474 ( .A(n338), .ZN(n242) );
  XNOR2_X1 U475 ( .A(n338), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U476 ( .A(n338), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U477 ( .A(n338), .B(n343), .ZN(n209) );
  XNOR2_X1 U478 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U479 ( .A(n292), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U480 ( .A(n338), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U481 ( .A(n36), .B(n3), .ZN(product[11]) );
  AOI21_X1 U482 ( .B1(n36), .B2(n332), .A(n304), .ZN(n31) );
  AOI21_X1 U483 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U484 ( .B1(n49), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U485 ( .A(n49), .ZN(n48) );
  OAI22_X1 U486 ( .A1(n340), .A2(n204), .B1(n203), .B2(n341), .ZN(n169) );
  OAI22_X1 U487 ( .A1(n340), .A2(n207), .B1(n206), .B2(n341), .ZN(n172) );
  OAI22_X1 U488 ( .A1(n340), .A2(n206), .B1(n205), .B2(n341), .ZN(n171) );
  OAI22_X1 U489 ( .A1(n340), .A2(n205), .B1(n204), .B2(n341), .ZN(n170) );
  OAI22_X1 U490 ( .A1(n340), .A2(n208), .B1(n207), .B2(n326), .ZN(n173) );
  OAI22_X1 U491 ( .A1(n340), .A2(n242), .B1(n210), .B2(n326), .ZN(n150) );
  OAI22_X1 U492 ( .A1(n234), .A2(n203), .B1(n296), .B2(n297), .ZN(n110) );
  XNOR2_X1 U493 ( .A(n336), .B(b[5]), .ZN(n213) );
  OAI22_X1 U494 ( .A1(n291), .A2(n234), .B1(n202), .B2(n341), .ZN(n142) );
  XNOR2_X1 U495 ( .A(n336), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U496 ( .A(n336), .B(b[4]), .ZN(n214) );
  INV_X1 U497 ( .A(n238), .ZN(n143) );
  OAI22_X1 U498 ( .A1(n340), .A2(n209), .B1(n208), .B2(n326), .ZN(n174) );
  XNOR2_X1 U499 ( .A(n336), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U500 ( .A(n343), .B(n336), .ZN(n218) );
  XNOR2_X1 U501 ( .A(n336), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U502 ( .A(n336), .B(b[2]), .ZN(n216) );
  INV_X1 U503 ( .A(n336), .ZN(n243) );
  XNOR2_X1 U504 ( .A(n336), .B(b[1]), .ZN(n217) );
  XOR2_X1 U505 ( .A(n247), .B(n146), .Z(n231) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n33, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86, n87,
         n88, n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n139, n140, n142, n143, n145, n146, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n240, n241, n242, n243, n244, n245, n246, n247,
         n255, n285, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n322), .B(n161), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n111), .B(n162), .CI(n156), .CO(n108), .S(n109) );
  FA_X1 U117 ( .A(n120), .B(n117), .CI(n115), .CO(n112), .S(n113) );
  FA_X1 U118 ( .A(n163), .B(n176), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U122 ( .A(n170), .B(n177), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n171), .B(n159), .CI(n178), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n181), .B(n174), .CO(n134), .S(n135) );
  BUF_X1 U249 ( .A(n244), .Z(n296) );
  BUF_X1 U250 ( .A(a[4]), .Z(n285) );
  BUF_X1 U251 ( .A(n237), .Z(n344) );
  BUF_X2 U252 ( .A(n347), .Z(n324) );
  INV_X1 U253 ( .A(n311), .ZN(n65) );
  AND2_X1 U254 ( .A1(n337), .A2(n80), .ZN(product[1]) );
  XNOR2_X1 U255 ( .A(n31), .B(n287), .ZN(product[12]) );
  AND2_X1 U256 ( .A1(n339), .A2(n30), .ZN(n287) );
  CLKBUF_X1 U257 ( .A(n332), .Z(n288) );
  CLKBUF_X1 U258 ( .A(n66), .Z(n289) );
  OAI21_X1 U259 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  INV_X1 U260 ( .A(n143), .ZN(n290) );
  CLKBUF_X1 U261 ( .A(b[7]), .Z(n291) );
  XNOR2_X1 U262 ( .A(n333), .B(b[7]), .ZN(n292) );
  INV_X1 U263 ( .A(n314), .ZN(n293) );
  BUF_X2 U264 ( .A(n238), .Z(n349) );
  CLKBUF_X1 U265 ( .A(n350), .Z(n294) );
  BUF_X2 U266 ( .A(n227), .Z(n350) );
  XOR2_X1 U267 ( .A(n241), .B(b[3]), .Z(n197) );
  XOR2_X1 U268 ( .A(n241), .B(b[6]), .Z(n194) );
  BUF_X2 U269 ( .A(n246), .Z(n295) );
  CLKBUF_X1 U270 ( .A(n246), .Z(n306) );
  AOI21_X1 U271 ( .B1(n326), .B2(n323), .A(n329), .ZN(n49) );
  BUF_X2 U272 ( .A(n247), .Z(n333) );
  XOR2_X1 U273 ( .A(n126), .B(n123), .Z(n297) );
  XOR2_X1 U274 ( .A(n121), .B(n297), .Z(n119) );
  NAND2_X1 U275 ( .A1(n121), .A2(n126), .ZN(n298) );
  NAND2_X1 U276 ( .A1(n121), .A2(n123), .ZN(n299) );
  NAND2_X1 U277 ( .A1(n126), .A2(n123), .ZN(n300) );
  NAND3_X1 U278 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n118) );
  XOR2_X1 U279 ( .A(n245), .B(n285), .Z(n301) );
  BUF_X1 U280 ( .A(n247), .Z(n342) );
  CLKBUF_X1 U281 ( .A(n336), .Z(n302) );
  CLKBUF_X1 U282 ( .A(n245), .Z(n303) );
  AOI21_X1 U283 ( .B1(n326), .B2(n58), .A(n329), .ZN(n304) );
  XOR2_X1 U284 ( .A(n342), .B(n146), .Z(n305) );
  OR2_X2 U285 ( .A1(n129), .A2(n132), .ZN(n338) );
  NAND2_X1 U286 ( .A1(n238), .A2(n230), .ZN(n307) );
  NAND2_X1 U287 ( .A1(n238), .A2(n230), .ZN(n234) );
  CLKBUF_X1 U288 ( .A(n232), .Z(n308) );
  XNOR2_X1 U289 ( .A(n245), .B(a[6]), .ZN(n309) );
  NOR2_X1 U290 ( .A1(n25), .A2(n20), .ZN(n310) );
  AND2_X2 U291 ( .A1(n129), .A2(n132), .ZN(n311) );
  NOR2_X2 U292 ( .A1(n103), .A2(n106), .ZN(n41) );
  BUF_X1 U293 ( .A(n237), .Z(n345) );
  CLKBUF_X1 U294 ( .A(n33), .Z(n312) );
  NAND2_X1 U295 ( .A1(n229), .A2(n344), .ZN(n313) );
  CLKBUF_X1 U296 ( .A(n245), .Z(n314) );
  XOR2_X1 U297 ( .A(n244), .B(a[6]), .Z(n315) );
  NAND2_X1 U298 ( .A1(n305), .A2(n255), .ZN(n316) );
  NAND2_X1 U299 ( .A1(n305), .A2(n255), .ZN(n317) );
  NAND2_X1 U300 ( .A1(n231), .A2(n255), .ZN(n235) );
  AOI21_X1 U301 ( .B1(n338), .B2(n66), .A(n311), .ZN(n318) );
  AOI21_X1 U302 ( .B1(n338), .B2(n289), .A(n311), .ZN(n319) );
  AOI21_X1 U303 ( .B1(n338), .B2(n66), .A(n311), .ZN(n61) );
  NAND2_X1 U304 ( .A1(n301), .A2(n344), .ZN(n320) );
  CLKBUF_X1 U305 ( .A(n53), .Z(n321) );
  OAI22_X1 U306 ( .A1(n234), .A2(n203), .B1(n349), .B2(n202), .ZN(n322) );
  OAI21_X1 U307 ( .B1(n59), .B2(n318), .A(n60), .ZN(n323) );
  XNOR2_X1 U308 ( .A(n245), .B(a[6]), .ZN(n347) );
  CLKBUF_X1 U309 ( .A(n302), .Z(n325) );
  NOR2_X1 U310 ( .A1(n335), .A2(n55), .ZN(n326) );
  CLKBUF_X1 U311 ( .A(n348), .Z(n327) );
  AOI21_X1 U312 ( .B1(n312), .B2(n339), .A(n28), .ZN(n328) );
  OAI21_X1 U313 ( .B1(n52), .B2(n56), .A(n53), .ZN(n329) );
  NOR2_X1 U314 ( .A1(n313), .A2(n198), .ZN(n330) );
  NOR2_X1 U315 ( .A1(n197), .A2(n345), .ZN(n331) );
  OR2_X1 U316 ( .A1(n330), .A2(n331), .ZN(n164) );
  OAI21_X1 U317 ( .B1(n49), .B2(n37), .A(n38), .ZN(n332) );
  AOI21_X1 U318 ( .B1(n50), .B2(n58), .A(n51), .ZN(n334) );
  NOR2_X1 U319 ( .A1(n113), .A2(n118), .ZN(n335) );
  NAND2_X1 U320 ( .A1(n236), .A2(n228), .ZN(n336) );
  OR2_X1 U321 ( .A1(n183), .A2(n151), .ZN(n337) );
  XNOR2_X1 U322 ( .A(n247), .B(a[2]), .ZN(n238) );
  INV_X1 U323 ( .A(n39), .ZN(n37) );
  INV_X1 U324 ( .A(n40), .ZN(n38) );
  NAND2_X1 U325 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U326 ( .A(n46), .ZN(n85) );
  INV_X1 U327 ( .A(n25), .ZN(n23) );
  INV_X1 U328 ( .A(n47), .ZN(n45) );
  INV_X1 U329 ( .A(n77), .ZN(n75) );
  NOR2_X1 U330 ( .A1(n113), .A2(n118), .ZN(n52) );
  NAND2_X1 U331 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U332 ( .A(n71), .ZN(n91) );
  NAND2_X1 U333 ( .A1(n107), .A2(n112), .ZN(n47) );
  AOI21_X1 U334 ( .B1(n33), .B2(n339), .A(n28), .ZN(n26) );
  INV_X1 U335 ( .A(n30), .ZN(n28) );
  INV_X1 U336 ( .A(n20), .ZN(n81) );
  XOR2_X1 U337 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U338 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U339 ( .A(n55), .ZN(n87) );
  XOR2_X1 U340 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U341 ( .A1(n84), .A2(n42), .ZN(n4) );
  XNOR2_X1 U342 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U343 ( .A1(n86), .A2(n321), .ZN(n6) );
  OAI21_X1 U344 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  INV_X1 U345 ( .A(n335), .ZN(n86) );
  XOR2_X1 U346 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U347 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U348 ( .A(n67), .ZN(n90) );
  XNOR2_X1 U349 ( .A(n9), .B(n289), .ZN(product[5]) );
  NAND2_X1 U350 ( .A1(n338), .A2(n65), .ZN(n9) );
  XNOR2_X1 U351 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U352 ( .A1(n340), .A2(n77), .ZN(n12) );
  NOR2_X1 U353 ( .A1(n25), .A2(n20), .ZN(n18) );
  INV_X1 U354 ( .A(n35), .ZN(n33) );
  NAND2_X1 U355 ( .A1(n113), .A2(n118), .ZN(n53) );
  INV_X1 U356 ( .A(n80), .ZN(n78) );
  XOR2_X1 U357 ( .A(n8), .B(n319), .Z(product[6]) );
  NAND2_X1 U358 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U359 ( .A(n59), .ZN(n88) );
  XNOR2_X1 U360 ( .A(n169), .B(n157), .ZN(n117) );
  NOR2_X1 U361 ( .A1(n96), .A2(n95), .ZN(n20) );
  NOR2_X1 U362 ( .A1(n124), .A2(n119), .ZN(n55) );
  INV_X1 U363 ( .A(n94), .ZN(n95) );
  OR2_X1 U364 ( .A1(n169), .A2(n157), .ZN(n116) );
  NAND2_X1 U365 ( .A1(n183), .A2(n151), .ZN(n80) );
  NAND2_X1 U366 ( .A1(n119), .A2(n124), .ZN(n56) );
  NOR2_X1 U367 ( .A1(n125), .A2(n128), .ZN(n59) );
  NOR2_X1 U368 ( .A1(n135), .A2(n150), .ZN(n71) );
  OR2_X1 U369 ( .A1(n98), .A2(n97), .ZN(n339) );
  NAND2_X1 U370 ( .A1(n125), .A2(n128), .ZN(n60) );
  OR2_X1 U371 ( .A1(n182), .A2(n175), .ZN(n340) );
  NAND2_X1 U372 ( .A1(n103), .A2(n106), .ZN(n42) );
  NAND2_X1 U373 ( .A1(n133), .A2(n134), .ZN(n68) );
  NAND2_X1 U374 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U375 ( .A1(n99), .A2(n102), .ZN(n341) );
  AND2_X1 U376 ( .A1(n294), .A2(n143), .ZN(n175) );
  INV_X1 U377 ( .A(n14), .ZN(product[15]) );
  OR2_X1 U378 ( .A1(n294), .A2(n242), .ZN(n210) );
  OAI22_X1 U379 ( .A1(n316), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OR2_X1 U380 ( .A1(n350), .A2(n243), .ZN(n219) );
  OAI22_X1 U381 ( .A1(n317), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  AND2_X1 U382 ( .A1(n350), .A2(n137), .ZN(n159) );
  OAI22_X1 U383 ( .A1(n316), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OR2_X1 U384 ( .A1(n294), .A2(n241), .ZN(n201) );
  OAI22_X1 U385 ( .A1(n316), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  AND2_X1 U386 ( .A1(n294), .A2(n140), .ZN(n167) );
  INV_X1 U387 ( .A(n139), .ZN(n160) );
  INV_X1 U388 ( .A(n100), .ZN(n101) );
  INV_X1 U389 ( .A(n136), .ZN(n152) );
  OR2_X1 U390 ( .A1(n350), .A2(n240), .ZN(n192) );
  INV_X1 U391 ( .A(n146), .ZN(n255) );
  NAND2_X1 U392 ( .A1(n309), .A2(n315), .ZN(n232) );
  AND2_X1 U393 ( .A1(n350), .A2(n146), .ZN(product[0]) );
  INV_X1 U394 ( .A(n145), .ZN(n176) );
  INV_X1 U395 ( .A(n142), .ZN(n168) );
  BUF_X1 U396 ( .A(n237), .Z(n343) );
  XNOR2_X1 U397 ( .A(n246), .B(a[4]), .ZN(n237) );
  NAND2_X1 U398 ( .A1(n135), .A2(n150), .ZN(n72) );
  OAI21_X1 U399 ( .B1(n41), .B2(n47), .A(n42), .ZN(n40) );
  INV_X1 U400 ( .A(n41), .ZN(n84) );
  NOR2_X1 U401 ( .A1(n46), .A2(n41), .ZN(n39) );
  XNOR2_X1 U402 ( .A(n22), .B(n346), .ZN(product[13]) );
  AND2_X1 U403 ( .A1(n81), .A2(n21), .ZN(n346) );
  OAI22_X1 U404 ( .A1(n317), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U405 ( .A1(n317), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  XNOR2_X1 U406 ( .A(n245), .B(a[6]), .ZN(n236) );
  XNOR2_X1 U407 ( .A(n296), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U408 ( .A(n296), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U409 ( .A(n296), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U410 ( .A(n350), .B(n244), .ZN(n191) );
  XNOR2_X1 U411 ( .A(n244), .B(b[1]), .ZN(n190) );
  INV_X1 U412 ( .A(n244), .ZN(n240) );
  XOR2_X1 U413 ( .A(n244), .B(a[6]), .Z(n228) );
  INV_X1 U414 ( .A(n110), .ZN(n111) );
  NOR2_X1 U415 ( .A1(n107), .A2(n112), .ZN(n46) );
  OAI22_X1 U416 ( .A1(n317), .A2(n212), .B1(n292), .B2(n255), .ZN(n177) );
  OAI22_X1 U417 ( .A1(n235), .A2(n292), .B1(n211), .B2(n255), .ZN(n145) );
  NAND2_X1 U418 ( .A1(n301), .A2(n344), .ZN(n348) );
  NAND2_X1 U419 ( .A1(n229), .A2(n345), .ZN(n233) );
  XNOR2_X1 U420 ( .A(n296), .B(b[6]), .ZN(n185) );
  INV_X1 U421 ( .A(n70), .ZN(n69) );
  NOR2_X1 U422 ( .A1(n133), .A2(n134), .ZN(n67) );
  XOR2_X1 U423 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U424 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  AOI21_X1 U425 ( .B1(n340), .B2(n78), .A(n75), .ZN(n73) );
  NAND2_X1 U426 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U427 ( .A1(n184), .A2(n325), .B1(n184), .B2(n324), .ZN(n136) );
  OAI22_X1 U428 ( .A1(n325), .A2(n185), .B1(n184), .B2(n324), .ZN(n94) );
  OAI22_X1 U429 ( .A1(n308), .A2(n188), .B1(n187), .B2(n324), .ZN(n155) );
  OAI22_X1 U430 ( .A1(n302), .A2(n187), .B1(n186), .B2(n324), .ZN(n154) );
  OAI22_X1 U431 ( .A1(n308), .A2(n186), .B1(n185), .B2(n324), .ZN(n153) );
  OAI22_X1 U432 ( .A1(n308), .A2(n190), .B1(n189), .B2(n324), .ZN(n157) );
  INV_X1 U433 ( .A(n347), .ZN(n137) );
  OAI22_X1 U434 ( .A1(n302), .A2(n189), .B1(n188), .B2(n324), .ZN(n156) );
  OAI22_X1 U435 ( .A1(n336), .A2(n240), .B1(n192), .B2(n347), .ZN(n148) );
  OAI22_X1 U436 ( .A1(n232), .A2(n191), .B1(n190), .B2(n347), .ZN(n158) );
  XNOR2_X1 U437 ( .A(n314), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U438 ( .A(n303), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U439 ( .A(n303), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U440 ( .A(n350), .B(n314), .ZN(n200) );
  XNOR2_X1 U441 ( .A(n303), .B(b[1]), .ZN(n199) );
  INV_X1 U442 ( .A(n245), .ZN(n241) );
  XOR2_X1 U443 ( .A(n245), .B(n285), .Z(n229) );
  INV_X1 U444 ( .A(n328), .ZN(n24) );
  OAI21_X1 U445 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U446 ( .A1(n98), .A2(n97), .ZN(n30) );
  OAI22_X1 U447 ( .A1(n327), .A2(n199), .B1(n198), .B2(n343), .ZN(n165) );
  OAI22_X1 U448 ( .A1(n320), .A2(n197), .B1(n343), .B2(n196), .ZN(n163) );
  INV_X1 U449 ( .A(n343), .ZN(n140) );
  OAI22_X1 U450 ( .A1(n320), .A2(n196), .B1(n195), .B2(n343), .ZN(n162) );
  OAI22_X1 U451 ( .A1(n348), .A2(n194), .B1(n193), .B2(n345), .ZN(n100) );
  XNOR2_X1 U452 ( .A(n295), .B(b[2]), .ZN(n207) );
  OAI22_X1 U453 ( .A1(n348), .A2(n293), .B1(n201), .B2(n343), .ZN(n149) );
  OAI22_X1 U454 ( .A1(n313), .A2(n200), .B1(n199), .B2(n343), .ZN(n166) );
  OAI22_X1 U455 ( .A1(n233), .A2(n195), .B1(n194), .B2(n343), .ZN(n161) );
  XNOR2_X1 U456 ( .A(n295), .B(b[5]), .ZN(n204) );
  XNOR2_X1 U457 ( .A(n295), .B(b[4]), .ZN(n205) );
  OAI22_X1 U458 ( .A1(n193), .A2(n327), .B1(n193), .B2(n343), .ZN(n139) );
  INV_X1 U459 ( .A(n295), .ZN(n242) );
  XNOR2_X1 U460 ( .A(n306), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U461 ( .A(n350), .B(n295), .ZN(n209) );
  XNOR2_X1 U462 ( .A(n295), .B(b[1]), .ZN(n208) );
  XOR2_X1 U463 ( .A(n246), .B(a[2]), .Z(n230) );
  XNOR2_X1 U464 ( .A(n296), .B(n291), .ZN(n184) );
  XNOR2_X1 U465 ( .A(n314), .B(n291), .ZN(n193) );
  XNOR2_X1 U466 ( .A(n306), .B(b[7]), .ZN(n202) );
  OAI21_X1 U467 ( .B1(n37), .B2(n49), .A(n38), .ZN(n36) );
  NAND2_X1 U468 ( .A1(n341), .A2(n35), .ZN(n3) );
  NAND2_X1 U469 ( .A1(n341), .A2(n339), .ZN(n25) );
  NAND2_X1 U470 ( .A1(n102), .A2(n99), .ZN(n35) );
  XNOR2_X1 U471 ( .A(n333), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U472 ( .A(n333), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U473 ( .A(n333), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U474 ( .A(n333), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U475 ( .A(n350), .B(n333), .ZN(n218) );
  XNOR2_X1 U476 ( .A(n333), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U477 ( .A(n333), .B(b[2]), .ZN(n216) );
  INV_X1 U478 ( .A(n333), .ZN(n243) );
  XOR2_X1 U479 ( .A(n146), .B(n342), .Z(n231) );
  XNOR2_X1 U480 ( .A(n48), .B(n5), .ZN(product[9]) );
  AOI21_X1 U481 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  INV_X1 U482 ( .A(n323), .ZN(n57) );
  OAI21_X1 U483 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  OAI21_X1 U484 ( .B1(n61), .B2(n59), .A(n60), .ZN(n58) );
  NOR2_X1 U485 ( .A1(n335), .A2(n55), .ZN(n50) );
  NAND2_X1 U486 ( .A1(n39), .A2(n310), .ZN(n16) );
  AOI21_X1 U487 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XNOR2_X1 U488 ( .A(n295), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U489 ( .A(n296), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U490 ( .A(n333), .B(b[3]), .ZN(n215) );
  OAI22_X1 U491 ( .A1(n316), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  XNOR2_X1 U492 ( .A(n288), .B(n3), .ZN(product[11]) );
  AOI21_X1 U493 ( .B1(n36), .B2(n341), .A(n312), .ZN(n31) );
  AOI21_X1 U494 ( .B1(n332), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U495 ( .B1(n334), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U496 ( .A(n304), .ZN(n48) );
  OAI22_X1 U497 ( .A1(n307), .A2(n204), .B1(n203), .B2(n290), .ZN(n169) );
  OAI22_X1 U498 ( .A1(n307), .A2(n207), .B1(n206), .B2(n290), .ZN(n172) );
  OAI22_X1 U499 ( .A1(n307), .A2(n206), .B1(n205), .B2(n349), .ZN(n171) );
  OAI22_X1 U500 ( .A1(n307), .A2(n205), .B1(n204), .B2(n349), .ZN(n170) );
  OAI22_X1 U501 ( .A1(n307), .A2(n208), .B1(n207), .B2(n349), .ZN(n173) );
  OAI22_X1 U502 ( .A1(n307), .A2(n242), .B1(n210), .B2(n290), .ZN(n150) );
  OAI22_X1 U503 ( .A1(n234), .A2(n203), .B1(n349), .B2(n202), .ZN(n110) );
  OAI22_X1 U504 ( .A1(n202), .A2(n234), .B1(n202), .B2(n349), .ZN(n142) );
  INV_X1 U505 ( .A(n349), .ZN(n143) );
  OAI22_X1 U506 ( .A1(n234), .A2(n209), .B1(n208), .B2(n349), .ZN(n174) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n24, n26, n28, n30, n31, n35, n36, n38, n39,
         n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n87, n88, n90, n91,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n139,
         n140, n142, n143, n145, n146, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n227, n230, n231, n232, n233, n234, n235, n238, n240, n241, n242,
         n243, n244, n245, n246, n247, n255, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n339, n340, n341, n342, n343, n344;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n328), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n156), .B(n162), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n164), .B(n177), .CI(n170), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  BUF_X1 U249 ( .A(n244), .Z(n299) );
  XNOR2_X1 U250 ( .A(n320), .B(b[5]), .ZN(n285) );
  BUF_X2 U251 ( .A(n245), .Z(n320) );
  AND2_X1 U252 ( .A1(n99), .A2(n102), .ZN(n317) );
  INV_X1 U253 ( .A(n317), .ZN(n35) );
  AND2_X1 U254 ( .A1(n335), .A2(n339), .ZN(n286) );
  OR2_X1 U255 ( .A1(n183), .A2(n151), .ZN(n287) );
  OR2_X1 U256 ( .A1(n46), .A2(n41), .ZN(n288) );
  NAND2_X1 U257 ( .A1(n307), .A2(n308), .ZN(n289) );
  OAI21_X1 U258 ( .B1(n52), .B2(n56), .A(n53), .ZN(n290) );
  OAI21_X1 U259 ( .B1(n294), .B2(n47), .A(n42), .ZN(n291) );
  CLKBUF_X1 U260 ( .A(n59), .Z(n292) );
  NOR2_X1 U261 ( .A1(n125), .A2(n128), .ZN(n59) );
  XOR2_X1 U262 ( .A(n246), .B(a[4]), .Z(n293) );
  NOR2_X1 U263 ( .A1(n103), .A2(n106), .ZN(n294) );
  INV_X1 U264 ( .A(n45), .ZN(n295) );
  CLKBUF_X1 U265 ( .A(n203), .Z(n296) );
  BUF_X2 U266 ( .A(n227), .Z(n297) );
  NAND2_X1 U267 ( .A1(n230), .A2(n238), .ZN(n298) );
  NAND2_X2 U268 ( .A1(n231), .A2(n255), .ZN(n235) );
  INV_X2 U269 ( .A(n146), .ZN(n255) );
  NOR2_X1 U270 ( .A1(n103), .A2(n106), .ZN(n41) );
  OR2_X2 U271 ( .A1(n330), .A2(n293), .ZN(n300) );
  OR2_X1 U272 ( .A1(n330), .A2(n331), .ZN(n233) );
  CLKBUF_X1 U273 ( .A(n246), .Z(n301) );
  NAND2_X1 U274 ( .A1(n333), .A2(n334), .ZN(n238) );
  NAND2_X2 U275 ( .A1(n333), .A2(n334), .ZN(n326) );
  OR2_X2 U276 ( .A1(n247), .A2(a[2]), .ZN(n334) );
  CLKBUF_X1 U277 ( .A(n246), .Z(n302) );
  XNOR2_X2 U278 ( .A(n246), .B(a[4]), .ZN(n343) );
  INV_X1 U279 ( .A(n243), .ZN(n303) );
  INV_X1 U280 ( .A(n243), .ZN(n304) );
  INV_X1 U281 ( .A(n243), .ZN(n344) );
  NAND2_X1 U282 ( .A1(a[2]), .A2(n306), .ZN(n307) );
  NAND2_X1 U283 ( .A1(n246), .A2(n305), .ZN(n308) );
  NAND2_X1 U284 ( .A1(n307), .A2(n308), .ZN(n230) );
  INV_X1 U285 ( .A(a[2]), .ZN(n305) );
  INV_X1 U286 ( .A(n246), .ZN(n306) );
  AOI21_X1 U287 ( .B1(n337), .B2(n66), .A(n63), .ZN(n309) );
  AOI21_X1 U288 ( .B1(n337), .B2(n66), .A(n63), .ZN(n310) );
  AOI21_X1 U289 ( .B1(n337), .B2(n66), .A(n63), .ZN(n61) );
  XNOR2_X1 U290 ( .A(n115), .B(n311), .ZN(n113) );
  XNOR2_X1 U291 ( .A(n120), .B(n117), .ZN(n311) );
  NAND2_X1 U292 ( .A1(n230), .A2(n238), .ZN(n312) );
  NAND2_X1 U293 ( .A1(n289), .A2(n238), .ZN(n234) );
  NAND2_X1 U294 ( .A1(n115), .A2(n120), .ZN(n313) );
  NAND2_X1 U295 ( .A1(n115), .A2(n117), .ZN(n314) );
  NAND2_X1 U296 ( .A1(n120), .A2(n117), .ZN(n315) );
  NAND3_X1 U297 ( .A1(n313), .A2(n314), .A3(n315), .ZN(n112) );
  CLKBUF_X1 U298 ( .A(n232), .Z(n316) );
  AND2_X1 U299 ( .A1(n335), .A2(n318), .ZN(n18) );
  AND2_X1 U300 ( .A1(n339), .A2(n81), .ZN(n318) );
  NOR2_X1 U301 ( .A1(n113), .A2(n118), .ZN(n319) );
  CLKBUF_X1 U302 ( .A(n246), .Z(n321) );
  XNOR2_X2 U303 ( .A(n245), .B(a[6]), .ZN(n341) );
  OR2_X2 U304 ( .A1(n323), .A2(n322), .ZN(n232) );
  XNOR2_X1 U305 ( .A(n244), .B(a[6]), .ZN(n322) );
  XOR2_X1 U306 ( .A(n245), .B(a[6]), .Z(n323) );
  OAI21_X1 U307 ( .B1(n61), .B2(n59), .A(n60), .ZN(n324) );
  OAI21_X1 U308 ( .B1(n59), .B2(n310), .A(n60), .ZN(n325) );
  CLKBUF_X1 U309 ( .A(n36), .Z(n327) );
  OAI22_X1 U310 ( .A1(n234), .A2(n203), .B1(n202), .B2(n326), .ZN(n328) );
  AOI21_X1 U311 ( .B1(n50), .B2(n325), .A(n51), .ZN(n329) );
  XNOR2_X1 U312 ( .A(n245), .B(a[4]), .ZN(n330) );
  XOR2_X1 U313 ( .A(n246), .B(a[4]), .Z(n331) );
  OAI22_X1 U314 ( .A1(n312), .A2(n203), .B1(n202), .B2(n326), .ZN(n110) );
  AOI21_X1 U315 ( .B1(n317), .B2(n339), .A(n28), .ZN(n332) );
  NAND2_X1 U316 ( .A1(n247), .A2(a[2]), .ZN(n333) );
  NAND2_X1 U317 ( .A1(n85), .A2(n295), .ZN(n5) );
  INV_X1 U318 ( .A(n46), .ZN(n85) );
  INV_X1 U319 ( .A(n47), .ZN(n45) );
  INV_X1 U320 ( .A(n77), .ZN(n75) );
  NOR2_X1 U321 ( .A1(n107), .A2(n112), .ZN(n46) );
  INV_X1 U322 ( .A(n30), .ZN(n28) );
  OAI21_X1 U323 ( .B1(n49), .B2(n288), .A(n38), .ZN(n36) );
  INV_X1 U324 ( .A(n291), .ZN(n38) );
  OAI21_X1 U325 ( .B1(n292), .B2(n309), .A(n60), .ZN(n58) );
  NAND2_X1 U326 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U327 ( .A(n20), .ZN(n81) );
  NAND2_X1 U328 ( .A1(n337), .A2(n65), .ZN(n9) );
  NAND2_X1 U329 ( .A1(n335), .A2(n35), .ZN(n3) );
  XOR2_X1 U330 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U331 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U332 ( .A(n41), .ZN(n84) );
  XOR2_X1 U333 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U334 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U335 ( .A(n55), .ZN(n87) );
  NAND2_X1 U336 ( .A1(n107), .A2(n112), .ZN(n47) );
  XNOR2_X1 U337 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U338 ( .A1(n336), .A2(n77), .ZN(n12) );
  NOR2_X1 U339 ( .A1(n46), .A2(n41), .ZN(n39) );
  INV_X1 U340 ( .A(n80), .ZN(n78) );
  NAND2_X1 U341 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U342 ( .A(n292), .ZN(n88) );
  INV_X1 U343 ( .A(n65), .ZN(n63) );
  AOI21_X1 U344 ( .B1(n50), .B2(n324), .A(n290), .ZN(n49) );
  OR2_X1 U345 ( .A1(n169), .A2(n157), .ZN(n116) );
  OAI21_X1 U346 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  NOR2_X1 U347 ( .A1(n119), .A2(n124), .ZN(n55) );
  INV_X1 U348 ( .A(n94), .ZN(n95) );
  NAND2_X1 U349 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U350 ( .A(n71), .ZN(n91) );
  XNOR2_X1 U351 ( .A(n169), .B(n157), .ZN(n117) );
  NOR2_X1 U352 ( .A1(n96), .A2(n95), .ZN(n20) );
  XOR2_X1 U353 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U354 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U355 ( .A(n67), .ZN(n90) );
  NAND2_X1 U356 ( .A1(n119), .A2(n124), .ZN(n56) );
  XNOR2_X1 U357 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U358 ( .A1(n342), .A2(n53), .ZN(n6) );
  OAI21_X1 U359 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  OR2_X1 U360 ( .A1(n99), .A2(n102), .ZN(n335) );
  NAND2_X1 U361 ( .A1(n125), .A2(n128), .ZN(n60) );
  INV_X1 U362 ( .A(n70), .ZN(n69) );
  NAND2_X1 U363 ( .A1(n96), .A2(n95), .ZN(n21) );
  NAND2_X1 U364 ( .A1(n103), .A2(n106), .ZN(n42) );
  OR2_X1 U365 ( .A1(n182), .A2(n175), .ZN(n336) );
  OR2_X1 U366 ( .A1(n129), .A2(n132), .ZN(n337) );
  AND2_X1 U367 ( .A1(n287), .A2(n80), .ZN(product[1]) );
  OR2_X1 U368 ( .A1(n98), .A2(n97), .ZN(n339) );
  INV_X1 U369 ( .A(n14), .ZN(product[15]) );
  AND2_X1 U370 ( .A1(n297), .A2(n140), .ZN(n167) );
  OAI22_X1 U371 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U372 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OR2_X1 U373 ( .A1(n297), .A2(n243), .ZN(n219) );
  OAI22_X1 U374 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OR2_X1 U375 ( .A1(n297), .A2(n241), .ZN(n201) );
  OAI22_X1 U376 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  NOR2_X1 U377 ( .A1(n133), .A2(n134), .ZN(n67) );
  INV_X1 U378 ( .A(n139), .ZN(n160) );
  INV_X1 U379 ( .A(n100), .ZN(n101) );
  INV_X1 U380 ( .A(n145), .ZN(n176) );
  OAI22_X1 U381 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  AND2_X1 U382 ( .A1(n297), .A2(n137), .ZN(n159) );
  OAI22_X1 U383 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  INV_X1 U384 ( .A(n136), .ZN(n152) );
  AND2_X1 U385 ( .A1(n297), .A2(n143), .ZN(n175) );
  NAND2_X1 U386 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U387 ( .A1(n297), .A2(n240), .ZN(n192) );
  OR2_X1 U388 ( .A1(n297), .A2(n242), .ZN(n210) );
  AND2_X1 U389 ( .A1(n297), .A2(n146), .ZN(product[0]) );
  NOR2_X1 U390 ( .A1(n135), .A2(n150), .ZN(n71) );
  INV_X1 U391 ( .A(n142), .ZN(n168) );
  CLKBUF_X1 U392 ( .A(n245), .Z(n340) );
  XNOR2_X1 U393 ( .A(n299), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U394 ( .A(n299), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U395 ( .A(n299), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U396 ( .A(n299), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U397 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U398 ( .A(n297), .B(n244), .ZN(n191) );
  INV_X1 U399 ( .A(n244), .ZN(n240) );
  AOI21_X1 U400 ( .B1(n336), .B2(n78), .A(n75), .ZN(n73) );
  OAI22_X1 U401 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OR2_X1 U402 ( .A1(n113), .A2(n118), .ZN(n342) );
  OAI22_X1 U403 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  INV_X1 U404 ( .A(n58), .ZN(n57) );
  XNOR2_X1 U405 ( .A(n9), .B(n66), .ZN(product[5]) );
  OAI22_X1 U406 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OAI21_X1 U407 ( .B1(n294), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U408 ( .A1(n129), .A2(n132), .ZN(n65) );
  XOR2_X1 U409 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U410 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  NAND2_X1 U411 ( .A1(n182), .A2(n175), .ZN(n77) );
  XNOR2_X1 U412 ( .A(n299), .B(b[2]), .ZN(n189) );
  NAND2_X1 U413 ( .A1(n339), .A2(n30), .ZN(n2) );
  AOI21_X1 U414 ( .B1(n317), .B2(n339), .A(n28), .ZN(n26) );
  NAND2_X1 U415 ( .A1(n98), .A2(n97), .ZN(n30) );
  OAI22_X1 U416 ( .A1(n300), .A2(n199), .B1(n198), .B2(n343), .ZN(n165) );
  OAI22_X1 U417 ( .A1(n300), .A2(n197), .B1(n196), .B2(n343), .ZN(n163) );
  OAI22_X1 U418 ( .A1(n233), .A2(n198), .B1(n197), .B2(n343), .ZN(n164) );
  OAI22_X1 U419 ( .A1(n300), .A2(n194), .B1(n193), .B2(n343), .ZN(n100) );
  OAI22_X1 U420 ( .A1(n300), .A2(n196), .B1(n195), .B2(n343), .ZN(n162) );
  INV_X1 U421 ( .A(n343), .ZN(n140) );
  OAI22_X1 U422 ( .A1(n233), .A2(n285), .B1(n194), .B2(n343), .ZN(n161) );
  OAI22_X1 U423 ( .A1(n300), .A2(n241), .B1(n201), .B2(n343), .ZN(n149) );
  OAI22_X1 U424 ( .A1(n233), .A2(n200), .B1(n199), .B2(n343), .ZN(n166) );
  OAI22_X1 U425 ( .A1(n193), .A2(n300), .B1(n193), .B2(n343), .ZN(n139) );
  INV_X1 U426 ( .A(n332), .ZN(n24) );
  OAI21_X1 U427 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  INV_X1 U428 ( .A(n110), .ZN(n111) );
  NOR2_X1 U429 ( .A1(n319), .A2(n55), .ZN(n50) );
  OAI22_X1 U430 ( .A1(n184), .A2(n316), .B1(n184), .B2(n341), .ZN(n136) );
  OAI21_X1 U431 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  NAND2_X1 U432 ( .A1(n113), .A2(n118), .ZN(n53) );
  NOR2_X1 U433 ( .A1(n113), .A2(n118), .ZN(n52) );
  OAI22_X1 U434 ( .A1(n316), .A2(n185), .B1(n184), .B2(n341), .ZN(n94) );
  OAI22_X1 U435 ( .A1(n316), .A2(n188), .B1(n187), .B2(n341), .ZN(n155) );
  OAI22_X1 U436 ( .A1(n232), .A2(n187), .B1(n186), .B2(n341), .ZN(n154) );
  OAI22_X1 U437 ( .A1(n232), .A2(n186), .B1(n185), .B2(n341), .ZN(n153) );
  OAI22_X1 U438 ( .A1(n232), .A2(n190), .B1(n189), .B2(n341), .ZN(n157) );
  INV_X1 U439 ( .A(n341), .ZN(n137) );
  OAI22_X1 U440 ( .A1(n232), .A2(n189), .B1(n188), .B2(n341), .ZN(n156) );
  OAI22_X1 U441 ( .A1(n232), .A2(n240), .B1(n192), .B2(n341), .ZN(n148) );
  OAI22_X1 U442 ( .A1(n232), .A2(n191), .B1(n190), .B2(n341), .ZN(n158) );
  XNOR2_X1 U443 ( .A(n340), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U444 ( .A(n340), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U445 ( .A(n320), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U446 ( .A(n340), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U447 ( .A(n320), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U448 ( .A(n297), .B(n320), .ZN(n200) );
  XNOR2_X1 U449 ( .A(n320), .B(b[6]), .ZN(n194) );
  INV_X1 U450 ( .A(n245), .ZN(n241) );
  NAND2_X1 U451 ( .A1(n39), .A2(n18), .ZN(n16) );
  AOI21_X1 U452 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XOR2_X1 U453 ( .A(n22), .B(n1), .Z(product[13]) );
  NAND2_X1 U454 ( .A1(n135), .A2(n150), .ZN(n72) );
  XOR2_X1 U455 ( .A(n31), .B(n2), .Z(product[12]) );
  XNOR2_X1 U456 ( .A(n321), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U457 ( .A(n321), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U458 ( .A(n302), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U459 ( .A(n302), .B(b[5]), .ZN(n204) );
  INV_X1 U460 ( .A(n321), .ZN(n242) );
  XNOR2_X1 U461 ( .A(n301), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U462 ( .A(n297), .B(n302), .ZN(n209) );
  XNOR2_X1 U463 ( .A(n246), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U464 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U465 ( .A(n8), .B(n309), .Z(product[6]) );
  AOI21_X1 U466 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  NAND2_X1 U467 ( .A1(n183), .A2(n151), .ZN(n80) );
  XNOR2_X1 U468 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U469 ( .A(n320), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U470 ( .A(n301), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U471 ( .A(n327), .B(n3), .ZN(product[11]) );
  AOI21_X1 U472 ( .B1(n36), .B2(n335), .A(n317), .ZN(n31) );
  AOI21_X1 U473 ( .B1(n36), .B2(n286), .A(n24), .ZN(n22) );
  OAI21_X1 U474 ( .B1(n329), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U475 ( .A(n49), .ZN(n48) );
  OAI22_X1 U476 ( .A1(n298), .A2(n204), .B1(n296), .B2(n326), .ZN(n169) );
  OAI22_X1 U477 ( .A1(n298), .A2(n207), .B1(n206), .B2(n326), .ZN(n172) );
  OAI22_X1 U478 ( .A1(n298), .A2(n206), .B1(n205), .B2(n326), .ZN(n171) );
  OAI22_X1 U479 ( .A1(n312), .A2(n205), .B1(n204), .B2(n326), .ZN(n170) );
  OAI22_X1 U480 ( .A1(n312), .A2(n208), .B1(n207), .B2(n326), .ZN(n173) );
  OAI22_X1 U481 ( .A1(n312), .A2(n242), .B1(n210), .B2(n326), .ZN(n150) );
  XNOR2_X1 U482 ( .A(n304), .B(b[5]), .ZN(n213) );
  OAI22_X1 U483 ( .A1(n202), .A2(n234), .B1(n202), .B2(n326), .ZN(n142) );
  XNOR2_X1 U484 ( .A(n304), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U485 ( .A(n303), .B(b[4]), .ZN(n214) );
  INV_X1 U486 ( .A(n326), .ZN(n143) );
  OAI22_X1 U487 ( .A1(n298), .A2(n209), .B1(n208), .B2(n326), .ZN(n174) );
  XNOR2_X1 U488 ( .A(n344), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U489 ( .A(n297), .B(n303), .ZN(n218) );
  XNOR2_X1 U490 ( .A(n344), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U491 ( .A(n304), .B(b[2]), .ZN(n216) );
  INV_X1 U492 ( .A(n247), .ZN(n243) );
  XNOR2_X1 U493 ( .A(n303), .B(b[1]), .ZN(n217) );
  XOR2_X1 U494 ( .A(n247), .B(n146), .Z(n231) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n63, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86, n87, n90,
         n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n131, n132, n133, n134, n135, n136, n137, n139, n140,
         n142, n143, n145, n146, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n227,
         n228, n231, n232, n233, n234, n235, n236, n238, n240, n241, n242,
         n243, n244, n245, n246, n247, n255, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n331, n332, n333, n334,
         n335, n336, n337, n338;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n323), .B(n161), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n111), .B(n162), .CI(n156), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n164), .B(n177), .CI(n170), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n286), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  AND2_X1 U249 ( .A1(n102), .A2(n99), .ZN(n303) );
  INV_X1 U250 ( .A(n303), .ZN(n35) );
  INV_X1 U251 ( .A(n242), .ZN(n285) );
  INV_X1 U252 ( .A(n242), .ZN(n336) );
  AND2_X1 U253 ( .A1(n292), .A2(n296), .ZN(n286) );
  OR2_X1 U254 ( .A1(n183), .A2(n151), .ZN(n287) );
  OR2_X2 U255 ( .A1(n308), .A2(n309), .ZN(n288) );
  OR2_X1 U256 ( .A1(n125), .A2(n128), .ZN(n289) );
  OR2_X1 U257 ( .A1(n297), .A2(n298), .ZN(n291) );
  CLKBUF_X1 U258 ( .A(n245), .Z(n290) );
  OAI22_X1 U259 ( .A1(n288), .A2(n241), .B1(n201), .B2(n335), .ZN(n292) );
  CLKBUF_X1 U260 ( .A(n246), .Z(n293) );
  BUF_X2 U261 ( .A(n238), .Z(n337) );
  CLKBUF_X1 U262 ( .A(n245), .Z(n294) );
  CLKBUF_X1 U263 ( .A(n66), .Z(n295) );
  OAI22_X1 U264 ( .A1(n288), .A2(n200), .B1(n199), .B2(n335), .ZN(n296) );
  XNOR2_X2 U265 ( .A(n246), .B(a[4]), .ZN(n335) );
  OR2_X2 U266 ( .A1(n297), .A2(n298), .ZN(n234) );
  XNOR2_X1 U267 ( .A(n246), .B(a[2]), .ZN(n297) );
  XOR2_X1 U268 ( .A(n247), .B(a[2]), .Z(n298) );
  XNOR2_X1 U269 ( .A(n31), .B(n299), .ZN(product[12]) );
  AND2_X1 U270 ( .A1(n301), .A2(n30), .ZN(n299) );
  XNOR2_X1 U271 ( .A(n22), .B(n300), .ZN(product[13]) );
  AND2_X1 U272 ( .A1(n81), .A2(n21), .ZN(n300) );
  CLKBUF_X1 U273 ( .A(n327), .Z(n301) );
  NOR2_X1 U274 ( .A1(n103), .A2(n106), .ZN(n302) );
  NOR2_X1 U275 ( .A1(n103), .A2(n106), .ZN(n41) );
  BUF_X2 U276 ( .A(n227), .Z(n338) );
  XNOR2_X1 U277 ( .A(n293), .B(b[6]), .ZN(n203) );
  XOR2_X1 U278 ( .A(n149), .B(n166), .Z(n131) );
  XNOR2_X1 U279 ( .A(n115), .B(n304), .ZN(n113) );
  XNOR2_X1 U280 ( .A(n120), .B(n117), .ZN(n304) );
  NOR2_X1 U281 ( .A1(n25), .A2(n20), .ZN(n305) );
  OAI21_X1 U282 ( .B1(n302), .B2(n47), .A(n42), .ZN(n306) );
  CLKBUF_X1 U283 ( .A(n314), .Z(n307) );
  XNOR2_X1 U284 ( .A(n293), .B(b[7]), .ZN(n202) );
  BUF_X1 U285 ( .A(n232), .Z(n332) );
  BUF_X2 U286 ( .A(n325), .Z(n334) );
  OR2_X2 U287 ( .A1(n308), .A2(n309), .ZN(n233) );
  XNOR2_X1 U288 ( .A(n245), .B(a[4]), .ZN(n308) );
  XOR2_X1 U289 ( .A(n246), .B(a[4]), .Z(n309) );
  CLKBUF_X1 U290 ( .A(b[5]), .Z(n310) );
  CLKBUF_X1 U291 ( .A(n247), .Z(n311) );
  AOI21_X1 U292 ( .B1(n328), .B2(n66), .A(n63), .ZN(n312) );
  AOI21_X1 U293 ( .B1(n328), .B2(n66), .A(n63), .ZN(n313) );
  OAI21_X1 U294 ( .B1(n59), .B2(n312), .A(n60), .ZN(n314) );
  INV_X1 U295 ( .A(n243), .ZN(n315) );
  NAND2_X1 U296 ( .A1(n115), .A2(n120), .ZN(n316) );
  NAND2_X1 U297 ( .A1(n115), .A2(n117), .ZN(n317) );
  NAND2_X1 U298 ( .A1(n120), .A2(n117), .ZN(n318) );
  NAND3_X1 U299 ( .A1(n316), .A2(n317), .A3(n318), .ZN(n112) );
  INV_X2 U300 ( .A(n240), .ZN(n319) );
  AOI21_X1 U301 ( .B1(n58), .B2(n50), .A(n51), .ZN(n320) );
  AOI21_X1 U302 ( .B1(n314), .B2(n50), .A(n51), .ZN(n49) );
  CLKBUF_X1 U303 ( .A(n36), .Z(n321) );
  AOI21_X1 U304 ( .B1(n303), .B2(n301), .A(n28), .ZN(n322) );
  OAI22_X1 U305 ( .A1(n234), .A2(n203), .B1(n202), .B2(n337), .ZN(n323) );
  NOR2_X1 U306 ( .A1(n113), .A2(n118), .ZN(n324) );
  XNOR2_X1 U307 ( .A(n245), .B(a[6]), .ZN(n325) );
  OAI21_X1 U308 ( .B1(n320), .B2(n37), .A(n38), .ZN(n36) );
  NOR2_X1 U309 ( .A1(n119), .A2(n124), .ZN(n55) );
  NOR2_X1 U310 ( .A1(n96), .A2(n95), .ZN(n20) );
  OR2_X1 U311 ( .A1(n99), .A2(n102), .ZN(n326) );
  INV_X1 U312 ( .A(n306), .ZN(n38) );
  INV_X1 U313 ( .A(n39), .ZN(n37) );
  NAND2_X1 U314 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U315 ( .A(n46), .ZN(n85) );
  INV_X1 U316 ( .A(n47), .ZN(n45) );
  INV_X1 U317 ( .A(n25), .ZN(n23) );
  INV_X1 U318 ( .A(n30), .ZN(n28) );
  NOR2_X1 U319 ( .A1(n107), .A2(n112), .ZN(n46) );
  INV_X1 U320 ( .A(n65), .ZN(n63) );
  NOR2_X1 U321 ( .A1(n113), .A2(n118), .ZN(n52) );
  OAI21_X1 U322 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  INV_X1 U323 ( .A(n71), .ZN(n91) );
  NAND2_X1 U324 ( .A1(n289), .A2(n60), .ZN(n8) );
  INV_X1 U325 ( .A(n20), .ZN(n81) );
  NAND2_X1 U326 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U327 ( .A(n302), .ZN(n84) );
  NAND2_X1 U328 ( .A1(n326), .A2(n35), .ZN(n3) );
  XOR2_X1 U329 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U330 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U331 ( .A(n67), .ZN(n90) );
  XOR2_X1 U332 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U333 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U334 ( .A(n55), .ZN(n87) );
  NAND2_X1 U335 ( .A1(n113), .A2(n118), .ZN(n53) );
  XNOR2_X1 U336 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U337 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U338 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  XNOR2_X1 U339 ( .A(n9), .B(n295), .ZN(product[5]) );
  NAND2_X1 U340 ( .A1(n328), .A2(n65), .ZN(n9) );
  XNOR2_X1 U341 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U342 ( .A1(n329), .A2(n77), .ZN(n12) );
  NOR2_X1 U343 ( .A1(n46), .A2(n41), .ZN(n39) );
  XNOR2_X1 U344 ( .A(n169), .B(n157), .ZN(n117) );
  NOR2_X1 U345 ( .A1(n133), .A2(n134), .ZN(n67) );
  OR2_X1 U346 ( .A1(n169), .A2(n157), .ZN(n116) );
  INV_X1 U347 ( .A(n94), .ZN(n95) );
  NAND2_X1 U348 ( .A1(n119), .A2(n124), .ZN(n56) );
  OR2_X1 U349 ( .A1(n98), .A2(n97), .ZN(n327) );
  NOR2_X1 U350 ( .A1(n125), .A2(n128), .ZN(n59) );
  NAND2_X1 U351 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U352 ( .A1(n129), .A2(n132), .ZN(n328) );
  NAND2_X1 U353 ( .A1(n125), .A2(n128), .ZN(n60) );
  NAND2_X1 U354 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U355 ( .A1(n175), .A2(n182), .ZN(n329) );
  NAND2_X1 U356 ( .A1(n103), .A2(n106), .ZN(n42) );
  AND2_X1 U357 ( .A1(n338), .A2(n143), .ZN(n175) );
  INV_X1 U358 ( .A(n14), .ZN(product[15]) );
  OR2_X1 U359 ( .A1(n338), .A2(n242), .ZN(n210) );
  AND2_X1 U360 ( .A1(n338), .A2(n140), .ZN(n167) );
  OAI22_X1 U361 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OR2_X1 U362 ( .A1(n338), .A2(n241), .ZN(n201) );
  INV_X1 U363 ( .A(n139), .ZN(n160) );
  INV_X1 U364 ( .A(n100), .ZN(n101) );
  AND2_X1 U365 ( .A1(n338), .A2(n137), .ZN(n159) );
  OAI22_X1 U366 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  INV_X1 U367 ( .A(n136), .ZN(n152) );
  OR2_X1 U368 ( .A1(n338), .A2(n240), .ZN(n192) );
  AND2_X1 U369 ( .A1(n287), .A2(n80), .ZN(product[1]) );
  OAI22_X1 U370 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OR2_X1 U371 ( .A1(n338), .A2(n243), .ZN(n219) );
  AND2_X1 U372 ( .A1(n338), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U373 ( .A(n245), .B(a[6]), .ZN(n236) );
  BUF_X1 U374 ( .A(n232), .Z(n331) );
  CLKBUF_X1 U375 ( .A(n232), .Z(n333) );
  NAND2_X1 U376 ( .A1(n228), .A2(n236), .ZN(n232) );
  INV_X1 U377 ( .A(n77), .ZN(n75) );
  INV_X1 U378 ( .A(n80), .ZN(n78) );
  XNOR2_X1 U379 ( .A(n338), .B(n244), .ZN(n191) );
  XNOR2_X1 U380 ( .A(n319), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U381 ( .A(n319), .B(n310), .ZN(n186) );
  XNOR2_X1 U382 ( .A(n319), .B(b[6]), .ZN(n185) );
  INV_X1 U383 ( .A(n244), .ZN(n240) );
  OAI22_X1 U384 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  INV_X1 U385 ( .A(n110), .ZN(n111) );
  INV_X1 U386 ( .A(n145), .ZN(n176) );
  INV_X1 U387 ( .A(n70), .ZN(n69) );
  XOR2_X1 U388 ( .A(n11), .B(n73), .Z(product[3]) );
  XOR2_X1 U389 ( .A(n244), .B(a[6]), .Z(n228) );
  OAI22_X1 U390 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U391 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U392 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U393 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  NAND2_X1 U394 ( .A1(n129), .A2(n132), .ZN(n65) );
  NOR2_X1 U395 ( .A1(n25), .A2(n20), .ZN(n18) );
  OAI21_X1 U396 ( .B1(n41), .B2(n47), .A(n42), .ZN(n40) );
  NOR2_X1 U397 ( .A1(n135), .A2(n150), .ZN(n71) );
  AOI21_X1 U398 ( .B1(n329), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U399 ( .A(n142), .ZN(n168) );
  NAND2_X1 U400 ( .A1(n107), .A2(n112), .ZN(n47) );
  AOI21_X1 U401 ( .B1(n303), .B2(n327), .A(n28), .ZN(n26) );
  NAND2_X1 U402 ( .A1(n326), .A2(n327), .ZN(n25) );
  NAND2_X1 U403 ( .A1(n98), .A2(n97), .ZN(n30) );
  NAND2_X1 U404 ( .A1(n91), .A2(n72), .ZN(n11) );
  OAI21_X1 U405 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  XNOR2_X1 U406 ( .A(n247), .B(a[2]), .ZN(n238) );
  NAND2_X2 U407 ( .A1(n231), .A2(n255), .ZN(n235) );
  NAND2_X1 U408 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U409 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OAI21_X1 U410 ( .B1(n59), .B2(n312), .A(n60), .ZN(n58) );
  INV_X1 U411 ( .A(n324), .ZN(n86) );
  NOR2_X1 U412 ( .A1(n324), .A2(n55), .ZN(n50) );
  OAI21_X1 U413 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  INV_X1 U414 ( .A(n322), .ZN(n24) );
  OAI21_X1 U415 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  OAI22_X1 U416 ( .A1(n288), .A2(n199), .B1(n198), .B2(n335), .ZN(n165) );
  OAI22_X1 U417 ( .A1(n288), .A2(n197), .B1(n196), .B2(n335), .ZN(n163) );
  OAI22_X1 U418 ( .A1(n233), .A2(n198), .B1(n197), .B2(n335), .ZN(n164) );
  INV_X1 U419 ( .A(n335), .ZN(n140) );
  OAI22_X1 U420 ( .A1(n288), .A2(n194), .B1(n193), .B2(n335), .ZN(n100) );
  OAI22_X1 U421 ( .A1(n193), .A2(n288), .B1(n193), .B2(n335), .ZN(n139) );
  OAI22_X1 U422 ( .A1(n233), .A2(n241), .B1(n201), .B2(n335), .ZN(n149) );
  OAI22_X1 U423 ( .A1(n233), .A2(n200), .B1(n199), .B2(n335), .ZN(n166) );
  OAI22_X1 U424 ( .A1(n288), .A2(n196), .B1(n195), .B2(n335), .ZN(n162) );
  XNOR2_X1 U425 ( .A(n336), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U426 ( .A(n336), .B(b[5]), .ZN(n204) );
  INV_X1 U427 ( .A(n246), .ZN(n242) );
  OAI22_X1 U428 ( .A1(n233), .A2(n195), .B1(n194), .B2(n335), .ZN(n161) );
  XNOR2_X1 U429 ( .A(n338), .B(n285), .ZN(n209) );
  OAI22_X1 U430 ( .A1(n184), .A2(n332), .B1(n184), .B2(n334), .ZN(n136) );
  OAI22_X1 U431 ( .A1(n333), .A2(n185), .B1(n184), .B2(n334), .ZN(n94) );
  OAI22_X1 U432 ( .A1(n332), .A2(n188), .B1(n187), .B2(n334), .ZN(n155) );
  OAI22_X1 U433 ( .A1(n332), .A2(n187), .B1(n186), .B2(n334), .ZN(n154) );
  INV_X1 U434 ( .A(n325), .ZN(n137) );
  OAI22_X1 U435 ( .A1(n333), .A2(n186), .B1(n185), .B2(n334), .ZN(n153) );
  OAI22_X1 U436 ( .A1(n333), .A2(n190), .B1(n189), .B2(n334), .ZN(n157) );
  OAI22_X1 U437 ( .A1(n332), .A2(n189), .B1(n188), .B2(n325), .ZN(n156) );
  OAI22_X1 U438 ( .A1(n331), .A2(n240), .B1(n192), .B2(n325), .ZN(n148) );
  OAI22_X1 U439 ( .A1(n331), .A2(n191), .B1(n190), .B2(n325), .ZN(n158) );
  XNOR2_X1 U440 ( .A(n338), .B(n294), .ZN(n200) );
  XNOR2_X1 U441 ( .A(n294), .B(b[4]), .ZN(n196) );
  INV_X1 U442 ( .A(n245), .ZN(n241) );
  XNOR2_X1 U443 ( .A(n290), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U444 ( .A(n245), .B(b[6]), .ZN(n194) );
  INV_X1 U445 ( .A(n307), .ZN(n57) );
  NAND2_X1 U446 ( .A1(n135), .A2(n150), .ZN(n72) );
  NAND2_X1 U447 ( .A1(n305), .A2(n39), .ZN(n16) );
  AOI21_X1 U448 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  XNOR2_X1 U449 ( .A(n319), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U450 ( .A(b[7]), .B(n294), .ZN(n193) );
  XOR2_X1 U451 ( .A(n8), .B(n313), .Z(product[6]) );
  NAND2_X1 U452 ( .A1(n183), .A2(n151), .ZN(n80) );
  XNOR2_X1 U453 ( .A(n315), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U454 ( .A(n311), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U455 ( .A(n315), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U456 ( .A(n311), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U457 ( .A(n338), .B(n315), .ZN(n218) );
  INV_X1 U458 ( .A(n247), .ZN(n243) );
  XOR2_X1 U459 ( .A(n247), .B(n146), .Z(n231) );
  XNOR2_X1 U460 ( .A(n285), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U461 ( .A(n319), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U462 ( .A(n290), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U463 ( .A(n311), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U464 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U465 ( .A(n43), .B(n4), .Z(product[10]) );
  AOI21_X1 U466 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  XNOR2_X1 U467 ( .A(n319), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U468 ( .A(n285), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U469 ( .A(n290), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U470 ( .A(n315), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U471 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U472 ( .A(n245), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U473 ( .A(n336), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U474 ( .A(b[1]), .B(n311), .ZN(n217) );
  XNOR2_X1 U475 ( .A(n321), .B(n3), .ZN(product[11]) );
  AOI21_X1 U476 ( .B1(n36), .B2(n326), .A(n303), .ZN(n31) );
  AOI21_X1 U477 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U478 ( .B1(n49), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U479 ( .A(n320), .ZN(n48) );
  OAI22_X1 U480 ( .A1(n291), .A2(n204), .B1(n203), .B2(n337), .ZN(n169) );
  OAI22_X1 U481 ( .A1(n291), .A2(n207), .B1(n206), .B2(n337), .ZN(n172) );
  OAI22_X1 U482 ( .A1(n291), .A2(n206), .B1(n205), .B2(n337), .ZN(n171) );
  OAI22_X1 U483 ( .A1(n291), .A2(n205), .B1(n204), .B2(n337), .ZN(n170) );
  OAI22_X1 U484 ( .A1(n291), .A2(n208), .B1(n207), .B2(n337), .ZN(n173) );
  OAI22_X1 U485 ( .A1(n291), .A2(n242), .B1(n210), .B2(n337), .ZN(n150) );
  OAI22_X1 U486 ( .A1(n234), .A2(n203), .B1(n202), .B2(n337), .ZN(n110) );
  OAI22_X1 U487 ( .A1(n202), .A2(n234), .B1(n202), .B2(n337), .ZN(n142) );
  INV_X1 U488 ( .A(n337), .ZN(n143) );
  OAI22_X1 U489 ( .A1(n291), .A2(n209), .B1(n208), .B2(n337), .ZN(n174) );
  INV_X2 U490 ( .A(n146), .ZN(n255) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_8_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  NOR2_X1 U106 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  OAI21_X1 U107 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  OR2_X1 U108 ( .A1(A[0]), .A2(B[0]), .ZN(n142) );
  CLKBUF_X1 U109 ( .A(n43), .Z(n143) );
  CLKBUF_X1 U110 ( .A(n35), .Z(n144) );
  CLKBUF_X1 U111 ( .A(n38), .Z(n145) );
  CLKBUF_X1 U112 ( .A(n27), .Z(n146) );
  AOI21_X1 U113 ( .B1(n144), .B2(n153), .A(n32), .ZN(n147) );
  AOI21_X1 U114 ( .B1(n67), .B2(n152), .A(n64), .ZN(n148) );
  AOI21_X1 U115 ( .B1(n59), .B2(n151), .A(n56), .ZN(n149) );
  XNOR2_X1 U116 ( .A(n16), .B(n150), .ZN(SUM[15]) );
  XOR2_X1 U117 ( .A(B[15]), .B(A[15]), .Z(n150) );
  INV_X1 U118 ( .A(n34), .ZN(n32) );
  AOI21_X1 U119 ( .B1(n51), .B2(n156), .A(n48), .ZN(n46) );
  INV_X1 U120 ( .A(n50), .ZN(n48) );
  AOI21_X1 U121 ( .B1(n67), .B2(n152), .A(n64), .ZN(n62) );
  INV_X1 U122 ( .A(n66), .ZN(n64) );
  AOI21_X1 U123 ( .B1(n59), .B2(n151), .A(n56), .ZN(n54) );
  INV_X1 U124 ( .A(n58), .ZN(n56) );
  OAI21_X1 U125 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  AOI21_X1 U126 ( .B1(n43), .B2(n155), .A(n40), .ZN(n38) );
  INV_X1 U127 ( .A(n42), .ZN(n40) );
  NAND2_X1 U128 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U129 ( .A(n36), .ZN(n78) );
  NAND2_X1 U130 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U131 ( .A(n28), .ZN(n76) );
  NAND2_X1 U132 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U133 ( .A(n52), .ZN(n82) );
  NAND2_X1 U134 ( .A1(n157), .A2(n26), .ZN(n3) );
  NAND2_X1 U135 ( .A1(n151), .A2(n58), .ZN(n11) );
  NAND2_X1 U136 ( .A1(n155), .A2(n42), .ZN(n7) );
  NAND2_X1 U137 ( .A1(n156), .A2(n50), .ZN(n9) );
  NAND2_X1 U138 ( .A1(n153), .A2(n34), .ZN(n5) );
  XOR2_X1 U139 ( .A(n148), .B(n12), .Z(SUM[3]) );
  NAND2_X1 U140 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U141 ( .A(n60), .ZN(n84) );
  XOR2_X1 U142 ( .A(n46), .B(n8), .Z(SUM[7]) );
  NAND2_X1 U143 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U144 ( .A(n44), .ZN(n80) );
  XOR2_X1 U145 ( .A(n14), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U146 ( .A1(n86), .A2(n69), .ZN(n14) );
  XNOR2_X1 U147 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  NAND2_X1 U148 ( .A1(n154), .A2(n20), .ZN(n2) );
  XNOR2_X1 U149 ( .A(n67), .B(n13), .ZN(SUM[2]) );
  NAND2_X1 U150 ( .A1(n152), .A2(n66), .ZN(n13) );
  INV_X1 U151 ( .A(n20), .ZN(n18) );
  NAND2_X1 U152 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  INV_X1 U153 ( .A(n26), .ZN(n24) );
  NOR2_X1 U154 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  OR2_X1 U155 ( .A1(A[4]), .A2(B[4]), .ZN(n151) );
  OR2_X1 U156 ( .A1(A[2]), .A2(B[2]), .ZN(n152) );
  NOR2_X1 U157 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U158 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U159 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NOR2_X1 U160 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NAND2_X1 U161 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U162 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U163 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U164 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U165 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  NAND2_X1 U166 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  OR2_X1 U167 ( .A1(A[10]), .A2(B[10]), .ZN(n153) );
  OR2_X1 U168 ( .A1(A[14]), .A2(B[14]), .ZN(n154) );
  OR2_X1 U169 ( .A1(A[8]), .A2(B[8]), .ZN(n155) );
  OR2_X1 U170 ( .A1(A[6]), .A2(B[6]), .ZN(n156) );
  OR2_X1 U171 ( .A1(A[12]), .A2(B[12]), .ZN(n157) );
  NAND2_X1 U172 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U173 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  NAND2_X1 U174 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U175 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  AND2_X1 U176 ( .A1(n142), .A2(n71), .ZN(SUM[0]) );
  NAND2_X1 U177 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  INV_X1 U178 ( .A(n68), .ZN(n86) );
  NAND2_X1 U179 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  XNOR2_X1 U180 ( .A(n143), .B(n7), .ZN(SUM[8]) );
  AOI21_X1 U181 ( .B1(n35), .B2(n153), .A(n32), .ZN(n30) );
  OAI21_X1 U182 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  OAI21_X1 U183 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XNOR2_X1 U184 ( .A(n51), .B(n9), .ZN(SUM[6]) );
  XOR2_X1 U185 ( .A(n147), .B(n4), .Z(SUM[11]) );
  XOR2_X1 U186 ( .A(n145), .B(n6), .Z(SUM[9]) );
  XNOR2_X1 U187 ( .A(n146), .B(n3), .ZN(SUM[12]) );
  OAI21_X1 U188 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  XNOR2_X1 U189 ( .A(n144), .B(n5), .ZN(SUM[10]) );
  XNOR2_X1 U190 ( .A(n59), .B(n11), .ZN(SUM[4]) );
  XOR2_X1 U191 ( .A(n149), .B(n10), .Z(SUM[5]) );
  INV_X1 U192 ( .A(n22), .ZN(n73) );
  OAI21_X1 U193 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X1 U194 ( .B1(n21), .B2(n154), .A(n18), .ZN(n16) );
  NAND2_X1 U195 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  AOI21_X1 U196 ( .B1(n27), .B2(n157), .A(n24), .ZN(n22) );
endmodule


module add_layer_WIDTH16_8 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_8_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n142, n143, n144, n145, n146, n147, n148, n150,
         n151, n152, n153, n154, n155, n156, n157;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  OR2_X1 U106 ( .A1(A[0]), .A2(B[0]), .ZN(n142) );
  CLKBUF_X1 U107 ( .A(n35), .Z(n143) );
  CLKBUF_X1 U108 ( .A(n62), .Z(n144) );
  CLKBUF_X1 U109 ( .A(n54), .Z(n145) );
  AOI21_X1 U110 ( .B1(n143), .B2(n153), .A(n32), .ZN(n146) );
  CLKBUF_X1 U111 ( .A(n38), .Z(n147) );
  XNOR2_X1 U112 ( .A(n16), .B(n148), .ZN(SUM[15]) );
  XOR2_X1 U113 ( .A(B[15]), .B(A[15]), .Z(n148) );
  AND2_X1 U114 ( .A1(n142), .A2(n71), .ZN(SUM[0]) );
  INV_X1 U115 ( .A(n42), .ZN(n40) );
  INV_X1 U116 ( .A(n34), .ZN(n32) );
  INV_X1 U117 ( .A(n66), .ZN(n64) );
  INV_X1 U118 ( .A(n58), .ZN(n56) );
  INV_X1 U119 ( .A(n50), .ZN(n48) );
  NAND2_X1 U120 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U121 ( .A(n44), .ZN(n80) );
  NAND2_X1 U122 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U123 ( .A(n28), .ZN(n76) );
  NAND2_X1 U124 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U125 ( .A(n60), .ZN(n84) );
  NAND2_X1 U126 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U127 ( .A(n52), .ZN(n82) );
  NAND2_X1 U128 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U129 ( .A(n36), .ZN(n78) );
  NAND2_X1 U130 ( .A1(n153), .A2(n34), .ZN(n5) );
  NAND2_X1 U131 ( .A1(n154), .A2(n26), .ZN(n3) );
  NAND2_X1 U132 ( .A1(n152), .A2(n58), .ZN(n11) );
  NAND2_X1 U133 ( .A1(n151), .A2(n50), .ZN(n9) );
  NAND2_X1 U134 ( .A1(n156), .A2(n66), .ZN(n13) );
  NAND2_X1 U135 ( .A1(n150), .A2(n42), .ZN(n7) );
  XOR2_X1 U136 ( .A(n14), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U137 ( .A1(n86), .A2(n69), .ZN(n14) );
  XNOR2_X1 U138 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  NAND2_X1 U139 ( .A1(n155), .A2(n20), .ZN(n2) );
  INV_X1 U140 ( .A(n20), .ZN(n18) );
  INV_X1 U141 ( .A(n22), .ZN(n73) );
  INV_X1 U142 ( .A(n26), .ZN(n24) );
  NOR2_X1 U143 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  NOR2_X1 U144 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U145 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U146 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NOR2_X1 U147 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NAND2_X1 U148 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  NAND2_X1 U149 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U150 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U151 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U152 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U153 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U154 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  OR2_X1 U155 ( .A1(A[8]), .A2(B[8]), .ZN(n150) );
  OR2_X1 U156 ( .A1(A[6]), .A2(B[6]), .ZN(n151) );
  OR2_X1 U157 ( .A1(A[4]), .A2(B[4]), .ZN(n152) );
  OR2_X1 U158 ( .A1(A[10]), .A2(B[10]), .ZN(n153) );
  OR2_X1 U159 ( .A1(A[12]), .A2(B[12]), .ZN(n154) );
  OR2_X1 U160 ( .A1(A[14]), .A2(B[14]), .ZN(n155) );
  OR2_X1 U161 ( .A1(A[2]), .A2(B[2]), .ZN(n156) );
  NAND2_X1 U162 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U163 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U164 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  NAND2_X1 U165 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U166 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  XNOR2_X1 U167 ( .A(n27), .B(n3), .ZN(SUM[12]) );
  CLKBUF_X1 U168 ( .A(n46), .Z(n157) );
  AOI21_X1 U169 ( .B1(n51), .B2(n151), .A(n48), .ZN(n46) );
  XNOR2_X1 U170 ( .A(n51), .B(n9), .ZN(SUM[6]) );
  OAI21_X1 U171 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  NAND2_X1 U172 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  XOR2_X1 U173 ( .A(n157), .B(n8), .Z(SUM[7]) );
  XOR2_X1 U174 ( .A(n145), .B(n10), .Z(SUM[5]) );
  INV_X1 U175 ( .A(n68), .ZN(n86) );
  AOI21_X1 U176 ( .B1(n59), .B2(n152), .A(n56), .ZN(n54) );
  NAND2_X1 U177 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  NOR2_X1 U178 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  XNOR2_X1 U179 ( .A(n59), .B(n11), .ZN(SUM[4]) );
  XOR2_X1 U180 ( .A(n147), .B(n6), .Z(SUM[9]) );
  OAI21_X1 U181 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  XNOR2_X1 U182 ( .A(n143), .B(n5), .ZN(SUM[10]) );
  XNOR2_X1 U183 ( .A(n67), .B(n13), .ZN(SUM[2]) );
  XNOR2_X1 U184 ( .A(n43), .B(n7), .ZN(SUM[8]) );
  XOR2_X1 U185 ( .A(n144), .B(n12), .Z(SUM[3]) );
  AOI21_X1 U186 ( .B1(n43), .B2(n150), .A(n40), .ZN(n38) );
  AOI21_X1 U187 ( .B1(n67), .B2(n156), .A(n64), .ZN(n62) );
  OAI21_X1 U188 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  OAI21_X1 U189 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  OAI21_X1 U190 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  AOI21_X1 U191 ( .B1(n35), .B2(n153), .A(n32), .ZN(n30) );
  AOI21_X1 U192 ( .B1(n27), .B2(n154), .A(n24), .ZN(n22) );
  OAI21_X1 U193 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U194 ( .B1(n21), .B2(n155), .A(n18), .ZN(n16) );
  XOR2_X1 U195 ( .A(n146), .B(n4), .Z(SUM[11]) );
endmodule


module add_layer_WIDTH16_7 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_7_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37,
         n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70,
         n71, n73, n75, n77, n79, n81, n82, n83, n84, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n71), .CO(n16), .S(SUM[14]) );
  AND2_X1 U104 ( .A1(n157), .A2(n70), .ZN(SUM[0]) );
  CLKBUF_X1 U105 ( .A(n41), .Z(n141) );
  CLKBUF_X1 U106 ( .A(n66), .Z(n142) );
  CLKBUF_X1 U107 ( .A(n30), .Z(n143) );
  AOI21_X1 U108 ( .B1(n58), .B2(n142), .A(n59), .ZN(n144) );
  AOI21_X1 U109 ( .B1(n143), .B2(n155), .A(n27), .ZN(n145) );
  CLKBUF_X1 U110 ( .A(n54), .Z(n146) );
  CLKBUF_X1 U111 ( .A(n38), .Z(n147) );
  AOI21_X1 U112 ( .B1(n54), .B2(n152), .A(n51), .ZN(n148) );
  AOI21_X1 U113 ( .B1(n38), .B2(n153), .A(n35), .ZN(n149) );
  NOR2_X1 U114 ( .A1(A[3]), .A2(B[3]), .ZN(n150) );
  INV_X1 U115 ( .A(n37), .ZN(n35) );
  INV_X1 U116 ( .A(n29), .ZN(n27) );
  INV_X1 U117 ( .A(n45), .ZN(n43) );
  AOI21_X1 U118 ( .B1(n146), .B2(n152), .A(n51), .ZN(n49) );
  INV_X1 U119 ( .A(n53), .ZN(n51) );
  AOI21_X1 U120 ( .B1(n58), .B2(n66), .A(n59), .ZN(n57) );
  NAND2_X1 U121 ( .A1(n73), .A2(n24), .ZN(n3) );
  INV_X1 U122 ( .A(n23), .ZN(n73) );
  NAND2_X1 U123 ( .A1(n155), .A2(n29), .ZN(n4) );
  NAND2_X1 U124 ( .A1(n156), .A2(n21), .ZN(n2) );
  NAND2_X1 U125 ( .A1(n77), .A2(n40), .ZN(n7) );
  INV_X1 U126 ( .A(n39), .ZN(n77) );
  NAND2_X1 U127 ( .A1(n75), .A2(n32), .ZN(n5) );
  INV_X1 U128 ( .A(n31), .ZN(n75) );
  XOR2_X1 U129 ( .A(n49), .B(n9), .Z(SUM[6]) );
  NAND2_X1 U130 ( .A1(n79), .A2(n48), .ZN(n9) );
  INV_X1 U131 ( .A(n47), .ZN(n79) );
  XOR2_X1 U132 ( .A(n65), .B(n13), .Z(SUM[2]) );
  NAND2_X1 U133 ( .A1(n83), .A2(n64), .ZN(n13) );
  INV_X1 U134 ( .A(n63), .ZN(n83) );
  NAND2_X1 U135 ( .A1(n153), .A2(n37), .ZN(n6) );
  NAND2_X1 U136 ( .A1(n154), .A2(n45), .ZN(n8) );
  XNOR2_X1 U137 ( .A(n62), .B(n12), .ZN(SUM[3]) );
  NAND2_X1 U138 ( .A1(n82), .A2(n61), .ZN(n12) );
  OAI21_X1 U139 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  NAND2_X1 U140 ( .A1(n84), .A2(n68), .ZN(n14) );
  NAND2_X1 U141 ( .A1(n152), .A2(n53), .ZN(n10) );
  NAND2_X1 U142 ( .A1(n81), .A2(n56), .ZN(n11) );
  INV_X1 U143 ( .A(n55), .ZN(n81) );
  NOR2_X1 U144 ( .A1(A[2]), .A2(B[2]), .ZN(n63) );
  NAND2_X1 U145 ( .A1(A[2]), .A2(B[2]), .ZN(n64) );
  XNOR2_X1 U146 ( .A(n16), .B(n151), .ZN(SUM[15]) );
  XNOR2_X1 U147 ( .A(B[15]), .B(A[15]), .ZN(n151) );
  NOR2_X1 U148 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  OR2_X1 U149 ( .A1(A[5]), .A2(B[5]), .ZN(n152) );
  NOR2_X1 U150 ( .A1(A[8]), .A2(B[8]), .ZN(n39) );
  NOR2_X1 U151 ( .A1(A[6]), .A2(B[6]), .ZN(n47) );
  NOR2_X1 U152 ( .A1(A[4]), .A2(B[4]), .ZN(n55) );
  NOR2_X1 U153 ( .A1(A[10]), .A2(B[10]), .ZN(n31) );
  NOR2_X1 U154 ( .A1(A[12]), .A2(B[12]), .ZN(n23) );
  INV_X1 U155 ( .A(n21), .ZN(n19) );
  NAND2_X1 U156 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U157 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U158 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U159 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U160 ( .A1(A[13]), .A2(B[13]), .ZN(n21) );
  OR2_X1 U161 ( .A1(A[9]), .A2(B[9]), .ZN(n153) );
  OR2_X1 U162 ( .A1(A[7]), .A2(B[7]), .ZN(n154) );
  OR2_X1 U163 ( .A1(A[11]), .A2(B[11]), .ZN(n155) );
  OR2_X1 U164 ( .A1(A[13]), .A2(B[13]), .ZN(n156) );
  NAND2_X1 U165 ( .A1(A[8]), .A2(B[8]), .ZN(n40) );
  NAND2_X1 U166 ( .A1(A[6]), .A2(B[6]), .ZN(n48) );
  NAND2_X1 U167 ( .A1(A[4]), .A2(B[4]), .ZN(n56) );
  NAND2_X1 U168 ( .A1(A[10]), .A2(B[10]), .ZN(n32) );
  NAND2_X1 U169 ( .A1(A[12]), .A2(B[12]), .ZN(n24) );
  NAND2_X1 U170 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  OR2_X1 U171 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  XOR2_X1 U172 ( .A(n14), .B(n70), .Z(SUM[1]) );
  XNOR2_X1 U173 ( .A(n146), .B(n10), .ZN(SUM[5]) );
  XNOR2_X1 U174 ( .A(n46), .B(n8), .ZN(SUM[7]) );
  OAI21_X1 U175 ( .B1(n148), .B2(n47), .A(n48), .ZN(n46) );
  XNOR2_X1 U176 ( .A(n147), .B(n6), .ZN(SUM[9]) );
  OAI21_X1 U177 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U178 ( .A1(A[0]), .A2(B[0]), .ZN(n70) );
  AOI21_X1 U179 ( .B1(n46), .B2(n154), .A(n43), .ZN(n41) );
  XOR2_X1 U180 ( .A(n141), .B(n7), .Z(SUM[8]) );
  INV_X1 U181 ( .A(n67), .ZN(n84) );
  INV_X1 U182 ( .A(n142), .ZN(n65) );
  NAND2_X1 U183 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  NOR2_X1 U184 ( .A1(A[1]), .A2(B[1]), .ZN(n67) );
  OAI21_X1 U185 ( .B1(n67), .B2(n70), .A(n68), .ZN(n66) );
  XOR2_X1 U186 ( .A(n33), .B(n5), .Z(SUM[10]) );
  AOI21_X1 U187 ( .B1(n147), .B2(n153), .A(n35), .ZN(n33) );
  XOR2_X1 U188 ( .A(n145), .B(n3), .Z(SUM[12]) );
  XOR2_X1 U189 ( .A(n144), .B(n11), .Z(SUM[4]) );
  INV_X1 U190 ( .A(n150), .ZN(n82) );
  OAI21_X1 U191 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  NOR2_X1 U192 ( .A1(n63), .A2(n150), .ZN(n58) );
  OAI21_X1 U193 ( .B1(n60), .B2(n64), .A(n61), .ZN(n59) );
  AOI21_X1 U194 ( .B1(n30), .B2(n155), .A(n27), .ZN(n25) );
  XNOR2_X1 U195 ( .A(n143), .B(n4), .ZN(SUM[11]) );
  OAI21_X1 U196 ( .B1(n149), .B2(n31), .A(n32), .ZN(n30) );
  INV_X1 U197 ( .A(n17), .ZN(n71) );
  XNOR2_X1 U198 ( .A(n22), .B(n2), .ZN(SUM[13]) );
  AOI21_X1 U199 ( .B1(n22), .B2(n156), .A(n19), .ZN(n17) );
  OAI21_X1 U200 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
endmodule


module add_layer_WIDTH16_2 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_2_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_2 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_2 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_2 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_8 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_7 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_2 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X2 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_2 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8 \genblk1[0].mult  ( .clk(clk), .ia(
        {\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7 \genblk1[1].mult  ( .clk(clk), .ia(
        {\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6 \genblk1[2].mult  ( .clk(clk), .ia(
        {\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5 \genblk1[3].mult  ( .clk(clk), .ia(
        {\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_2 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86, n87,
         n88, n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n139, n140, n142, n143, n145, n146, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n240, n241, n242, n243, n244, n245, n246, n247,
         n255, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n334, n335, n336, n337, n338, n339,
         n340, n341, n342;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n302), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U115 ( .A(n156), .B(n162), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n170), .B(n177), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n166), .B(n149), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  BUF_X4 U249 ( .A(n246), .Z(n340) );
  AND2_X1 U250 ( .A1(n99), .A2(n102), .ZN(n314) );
  BUF_X2 U251 ( .A(n238), .Z(n336) );
  XNOR2_X1 U252 ( .A(n169), .B(n157), .ZN(n117) );
  OAI22_X1 U253 ( .A1(n321), .A2(n187), .B1(n186), .B2(n338), .ZN(n154) );
  INV_X1 U254 ( .A(n314), .ZN(n35) );
  OR2_X1 U255 ( .A1(n183), .A2(n151), .ZN(n285) );
  XOR2_X1 U256 ( .A(n241), .B(b[5]), .Z(n195) );
  BUF_X2 U257 ( .A(n237), .Z(n335) );
  INV_X1 U258 ( .A(n240), .ZN(n286) );
  INV_X1 U259 ( .A(n87), .ZN(n287) );
  OAI21_X1 U260 ( .B1(n297), .B2(n47), .A(n42), .ZN(n288) );
  NAND2_X1 U261 ( .A1(n231), .A2(n255), .ZN(n289) );
  XNOR2_X1 U262 ( .A(n246), .B(a[4]), .ZN(n290) );
  CLKBUF_X1 U263 ( .A(n342), .Z(n291) );
  CLKBUF_X1 U264 ( .A(n36), .Z(n326) );
  INV_X1 U265 ( .A(n241), .ZN(n292) );
  INV_X1 U266 ( .A(n312), .ZN(n313) );
  XNOR2_X1 U267 ( .A(n340), .B(b[7]), .ZN(n293) );
  XNOR2_X1 U268 ( .A(n115), .B(n294), .ZN(n113) );
  XNOR2_X1 U269 ( .A(n120), .B(n117), .ZN(n294) );
  CLKBUF_X1 U270 ( .A(n341), .Z(n295) );
  CLKBUF_X1 U271 ( .A(n58), .Z(n296) );
  NOR2_X1 U272 ( .A1(n103), .A2(n106), .ZN(n297) );
  BUF_X2 U273 ( .A(n247), .Z(n319) );
  CLKBUF_X1 U274 ( .A(n247), .Z(n310) );
  XNOR2_X1 U275 ( .A(n109), .B(n298), .ZN(n107) );
  XNOR2_X1 U276 ( .A(n114), .B(n116), .ZN(n298) );
  NAND2_X1 U277 ( .A1(n115), .A2(n120), .ZN(n299) );
  NAND2_X1 U278 ( .A1(n115), .A2(n117), .ZN(n300) );
  NAND2_X1 U279 ( .A1(n120), .A2(n117), .ZN(n301) );
  NAND3_X1 U280 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n112) );
  OAI22_X1 U281 ( .A1(n341), .A2(n203), .B1(n293), .B2(n336), .ZN(n302) );
  XNOR2_X1 U282 ( .A(n31), .B(n303), .ZN(product[12]) );
  AND2_X1 U283 ( .A1(n330), .A2(n30), .ZN(n303) );
  XNOR2_X1 U284 ( .A(n22), .B(n304), .ZN(product[13]) );
  AND2_X1 U285 ( .A1(n81), .A2(n21), .ZN(n304) );
  AOI21_X1 U286 ( .B1(n329), .B2(n66), .A(n63), .ZN(n305) );
  NAND2_X1 U287 ( .A1(n229), .A2(n290), .ZN(n306) );
  AOI21_X1 U288 ( .B1(n329), .B2(n66), .A(n63), .ZN(n61) );
  NAND2_X1 U289 ( .A1(n290), .A2(n229), .ZN(n233) );
  BUF_X2 U290 ( .A(n227), .Z(n342) );
  OAI21_X2 U291 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  NAND2_X1 U292 ( .A1(n109), .A2(n114), .ZN(n307) );
  NAND2_X1 U293 ( .A1(n109), .A2(n116), .ZN(n308) );
  NAND2_X1 U294 ( .A1(n114), .A2(n116), .ZN(n309) );
  NAND3_X1 U295 ( .A1(n307), .A2(n308), .A3(n309), .ZN(n106) );
  NOR2_X1 U296 ( .A1(n103), .A2(n106), .ZN(n41) );
  NOR2_X1 U297 ( .A1(n113), .A2(n118), .ZN(n311) );
  INV_X1 U298 ( .A(n245), .ZN(n312) );
  NOR2_X1 U299 ( .A1(n113), .A2(n118), .ZN(n52) );
  XOR2_X1 U300 ( .A(n101), .B(n154), .Z(n315) );
  XOR2_X1 U301 ( .A(n104), .B(n315), .Z(n99) );
  NAND2_X1 U302 ( .A1(n104), .A2(n101), .ZN(n316) );
  NAND2_X1 U303 ( .A1(n104), .A2(n154), .ZN(n317) );
  NAND2_X1 U304 ( .A1(n101), .A2(n154), .ZN(n318) );
  NAND3_X1 U305 ( .A1(n316), .A2(n317), .A3(n318), .ZN(n98) );
  OR2_X2 U306 ( .A1(n98), .A2(n97), .ZN(n330) );
  NAND2_X1 U307 ( .A1(n228), .A2(n327), .ZN(n320) );
  NAND2_X1 U308 ( .A1(n228), .A2(n327), .ZN(n321) );
  NAND2_X1 U309 ( .A1(n228), .A2(n327), .ZN(n232) );
  NAND2_X1 U310 ( .A1(n244), .A2(n323), .ZN(n324) );
  NAND2_X1 U311 ( .A1(n322), .A2(a[6]), .ZN(n325) );
  NAND2_X1 U312 ( .A1(n324), .A2(n325), .ZN(n228) );
  INV_X1 U313 ( .A(n244), .ZN(n322) );
  INV_X1 U314 ( .A(a[6]), .ZN(n323) );
  XNOR2_X1 U315 ( .A(n245), .B(a[6]), .ZN(n327) );
  AOI21_X1 U316 ( .B1(n58), .B2(n50), .A(n51), .ZN(n328) );
  XNOR2_X1 U317 ( .A(n326), .B(n3), .ZN(product[11]) );
  NOR2_X1 U318 ( .A1(n119), .A2(n124), .ZN(n55) );
  NAND2_X1 U319 ( .A1(n119), .A2(n124), .ZN(n56) );
  OR2_X1 U320 ( .A1(n129), .A2(n132), .ZN(n329) );
  INV_X1 U321 ( .A(n288), .ZN(n38) );
  INV_X1 U322 ( .A(n39), .ZN(n37) );
  XNOR2_X1 U323 ( .A(n48), .B(n5), .ZN(product[9]) );
  NAND2_X1 U324 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U325 ( .A(n46), .ZN(n85) );
  INV_X1 U326 ( .A(n47), .ZN(n45) );
  INV_X1 U327 ( .A(n65), .ZN(n63) );
  INV_X1 U328 ( .A(n77), .ZN(n75) );
  NOR2_X1 U329 ( .A1(n112), .A2(n107), .ZN(n46) );
  OAI21_X1 U330 ( .B1(n297), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U331 ( .A1(n107), .A2(n112), .ZN(n47) );
  NAND2_X1 U332 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U333 ( .A(n71), .ZN(n91) );
  NAND2_X1 U334 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U335 ( .A(n59), .ZN(n88) );
  INV_X1 U336 ( .A(n20), .ZN(n81) );
  NAND2_X1 U337 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U338 ( .A(n41), .ZN(n84) );
  NAND2_X1 U339 ( .A1(n329), .A2(n65), .ZN(n9) );
  XOR2_X1 U340 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U341 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U342 ( .A(n67), .ZN(n90) );
  XOR2_X1 U343 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U344 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U345 ( .A(n55), .ZN(n87) );
  XNOR2_X1 U346 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U347 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U348 ( .B1(n57), .B2(n287), .A(n56), .ZN(n54) );
  NOR2_X1 U349 ( .A1(n46), .A2(n41), .ZN(n39) );
  XNOR2_X1 U350 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U351 ( .A1(n332), .A2(n77), .ZN(n12) );
  INV_X1 U352 ( .A(n30), .ZN(n28) );
  NOR2_X1 U353 ( .A1(n96), .A2(n95), .ZN(n20) );
  OR2_X1 U354 ( .A1(n99), .A2(n102), .ZN(n331) );
  NOR2_X1 U355 ( .A1(n125), .A2(n128), .ZN(n59) );
  NOR2_X1 U356 ( .A1(n133), .A2(n134), .ZN(n67) );
  NOR2_X1 U357 ( .A1(n135), .A2(n150), .ZN(n71) );
  INV_X1 U358 ( .A(n80), .ZN(n78) );
  NAND2_X1 U359 ( .A1(n125), .A2(n128), .ZN(n60) );
  NAND2_X1 U360 ( .A1(n103), .A2(n106), .ZN(n42) );
  NAND2_X1 U361 ( .A1(n133), .A2(n134), .ZN(n68) );
  NAND2_X1 U362 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U363 ( .A1(n182), .A2(n175), .ZN(n332) );
  AND2_X1 U364 ( .A1(n342), .A2(n143), .ZN(n175) );
  INV_X1 U365 ( .A(n14), .ZN(product[15]) );
  OR2_X1 U366 ( .A1(n342), .A2(n242), .ZN(n210) );
  INV_X1 U367 ( .A(n340), .ZN(n242) );
  XNOR2_X1 U368 ( .A(n342), .B(n340), .ZN(n209) );
  AND2_X1 U369 ( .A1(n291), .A2(n140), .ZN(n167) );
  INV_X1 U370 ( .A(n110), .ZN(n111) );
  INV_X1 U371 ( .A(n145), .ZN(n176) );
  CLKBUF_X1 U372 ( .A(n237), .Z(n334) );
  OR2_X1 U373 ( .A1(n342), .A2(n240), .ZN(n192) );
  AND2_X1 U374 ( .A1(n285), .A2(n80), .ZN(product[1]) );
  OR2_X1 U375 ( .A1(n342), .A2(n243), .ZN(n219) );
  XNOR2_X1 U376 ( .A(n340), .B(b[5]), .ZN(n204) );
  XNOR2_X1 U377 ( .A(n340), .B(b[4]), .ZN(n205) );
  NAND2_X1 U378 ( .A1(n231), .A2(n255), .ZN(n235) );
  XNOR2_X1 U379 ( .A(n340), .B(b[7]), .ZN(n202) );
  XOR2_X1 U380 ( .A(n246), .B(a[2]), .Z(n230) );
  XNOR2_X1 U381 ( .A(n340), .B(b[3]), .ZN(n206) );
  AND2_X1 U382 ( .A1(n291), .A2(n146), .ZN(product[0]) );
  NAND2_X1 U383 ( .A1(n135), .A2(n150), .ZN(n72) );
  BUF_X1 U384 ( .A(n236), .Z(n337) );
  XNOR2_X1 U385 ( .A(n246), .B(a[4]), .ZN(n237) );
  XNOR2_X1 U386 ( .A(n286), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U387 ( .A(n286), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U388 ( .A(n244), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U389 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U390 ( .A(n342), .B(n244), .ZN(n191) );
  INV_X1 U391 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U392 ( .A(n247), .B(a[2]), .ZN(n238) );
  BUF_X2 U393 ( .A(n236), .Z(n338) );
  XNOR2_X1 U394 ( .A(n245), .B(a[6]), .ZN(n236) );
  NAND2_X1 U395 ( .A1(n331), .A2(n35), .ZN(n3) );
  INV_X1 U396 ( .A(n25), .ZN(n23) );
  OR2_X1 U397 ( .A1(n342), .A2(n241), .ZN(n201) );
  INV_X1 U398 ( .A(n136), .ZN(n152) );
  INV_X1 U399 ( .A(n94), .ZN(n95) );
  OR2_X1 U400 ( .A1(n169), .A2(n157), .ZN(n116) );
  AND2_X1 U401 ( .A1(n342), .A2(n137), .ZN(n159) );
  INV_X1 U402 ( .A(n100), .ZN(n101) );
  INV_X1 U403 ( .A(n139), .ZN(n160) );
  AOI21_X1 U404 ( .B1(n314), .B2(n330), .A(n28), .ZN(n339) );
  OAI21_X1 U405 ( .B1(n49), .B2(n37), .A(n38), .ZN(n36) );
  OAI22_X1 U406 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U407 ( .A1(n289), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U408 ( .A1(n289), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U409 ( .A1(n289), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OAI22_X1 U410 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U411 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  OAI22_X1 U412 ( .A1(n211), .A2(n289), .B1(n211), .B2(n255), .ZN(n145) );
  INV_X1 U413 ( .A(n339), .ZN(n24) );
  NAND2_X1 U414 ( .A1(n98), .A2(n97), .ZN(n30) );
  XOR2_X1 U415 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U416 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  AOI21_X1 U417 ( .B1(n332), .B2(n78), .A(n75), .ZN(n73) );
  NAND2_X1 U418 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U419 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  XNOR2_X1 U420 ( .A(n286), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U421 ( .A(n340), .B(b[6]), .ZN(n203) );
  NAND2_X1 U422 ( .A1(n230), .A2(n238), .ZN(n341) );
  NAND2_X1 U423 ( .A1(n238), .A2(n230), .ZN(n234) );
  INV_X1 U424 ( .A(n70), .ZN(n69) );
  XNOR2_X1 U425 ( .A(n340), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U426 ( .A(n244), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U427 ( .A(n9), .B(n66), .ZN(product[5]) );
  NAND2_X1 U428 ( .A1(n183), .A2(n151), .ZN(n80) );
  XOR2_X1 U429 ( .A(n245), .B(a[4]), .Z(n229) );
  INV_X1 U430 ( .A(n245), .ZN(n241) );
  XNOR2_X1 U431 ( .A(n292), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U432 ( .A(n313), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U433 ( .A(n292), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U434 ( .A(n313), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U435 ( .A(n292), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U436 ( .A(n342), .B(n313), .ZN(n200) );
  INV_X1 U437 ( .A(n142), .ZN(n168) );
  INV_X1 U438 ( .A(n296), .ZN(n57) );
  OAI21_X1 U439 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  XOR2_X1 U440 ( .A(n8), .B(n305), .Z(product[6]) );
  OAI22_X1 U441 ( .A1(n184), .A2(n320), .B1(n184), .B2(n337), .ZN(n136) );
  OAI22_X1 U442 ( .A1(n321), .A2(n185), .B1(n184), .B2(n338), .ZN(n94) );
  OAI22_X1 U443 ( .A1(n320), .A2(n188), .B1(n187), .B2(n337), .ZN(n155) );
  OAI22_X1 U444 ( .A1(n321), .A2(n190), .B1(n189), .B2(n338), .ZN(n157) );
  OAI22_X1 U445 ( .A1(n320), .A2(n186), .B1(n185), .B2(n337), .ZN(n153) );
  OAI22_X1 U446 ( .A1(n320), .A2(n189), .B1(n188), .B2(n337), .ZN(n156) );
  OAI22_X1 U447 ( .A1(n232), .A2(n240), .B1(n192), .B2(n337), .ZN(n148) );
  OAI22_X1 U448 ( .A1(n191), .A2(n232), .B1(n190), .B2(n338), .ZN(n158) );
  INV_X1 U449 ( .A(n338), .ZN(n137) );
  NAND2_X1 U450 ( .A1(n113), .A2(n118), .ZN(n53) );
  OAI21_X1 U451 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  AOI21_X1 U452 ( .B1(n314), .B2(n330), .A(n28), .ZN(n26) );
  OAI22_X1 U453 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  XOR2_X1 U454 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U455 ( .A1(n129), .A2(n132), .ZN(n65) );
  OAI22_X1 U456 ( .A1(n306), .A2(n199), .B1(n198), .B2(n334), .ZN(n165) );
  OAI22_X1 U457 ( .A1(n306), .A2(n197), .B1(n196), .B2(n335), .ZN(n163) );
  OAI22_X1 U458 ( .A1(n306), .A2(n198), .B1(n197), .B2(n334), .ZN(n164) );
  OAI22_X1 U459 ( .A1(n233), .A2(n194), .B1(n193), .B2(n334), .ZN(n100) );
  OAI22_X1 U460 ( .A1(n193), .A2(n306), .B1(n193), .B2(n335), .ZN(n139) );
  OAI22_X1 U461 ( .A1(n306), .A2(n196), .B1(n195), .B2(n334), .ZN(n162) );
  OAI22_X1 U462 ( .A1(n233), .A2(n195), .B1(n194), .B2(n334), .ZN(n161) );
  INV_X1 U463 ( .A(n335), .ZN(n140) );
  OAI22_X1 U464 ( .A1(n233), .A2(n241), .B1(n201), .B2(n335), .ZN(n149) );
  OAI22_X1 U465 ( .A1(n233), .A2(n200), .B1(n199), .B2(n335), .ZN(n166) );
  AOI21_X1 U466 ( .B1(n58), .B2(n50), .A(n51), .ZN(n49) );
  AOI21_X1 U467 ( .B1(n18), .B2(n40), .A(n19), .ZN(n17) );
  OAI21_X1 U468 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  NOR2_X1 U469 ( .A1(n311), .A2(n55), .ZN(n50) );
  INV_X1 U470 ( .A(n311), .ZN(n86) );
  NOR2_X1 U471 ( .A1(n25), .A2(n20), .ZN(n18) );
  NAND2_X1 U472 ( .A1(n331), .A2(n330), .ZN(n25) );
  NAND2_X1 U473 ( .A1(n39), .A2(n18), .ZN(n16) );
  AOI21_X1 U474 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  XNOR2_X1 U475 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U476 ( .A(n245), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U477 ( .A(n340), .B(b[1]), .ZN(n208) );
  AOI21_X1 U478 ( .B1(n36), .B2(n331), .A(n314), .ZN(n31) );
  AOI21_X1 U479 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U480 ( .B1(n328), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U481 ( .A(n49), .ZN(n48) );
  OAI22_X1 U482 ( .A1(n234), .A2(n204), .B1(n203), .B2(n336), .ZN(n169) );
  OAI22_X1 U483 ( .A1(n295), .A2(n207), .B1(n206), .B2(n336), .ZN(n172) );
  OAI22_X1 U484 ( .A1(n341), .A2(n206), .B1(n205), .B2(n336), .ZN(n171) );
  OAI22_X1 U485 ( .A1(n234), .A2(n205), .B1(n204), .B2(n336), .ZN(n170) );
  OAI22_X1 U486 ( .A1(n234), .A2(n208), .B1(n207), .B2(n336), .ZN(n173) );
  OAI22_X1 U487 ( .A1(n295), .A2(n242), .B1(n210), .B2(n336), .ZN(n150) );
  OAI22_X1 U488 ( .A1(n341), .A2(n203), .B1(n202), .B2(n336), .ZN(n110) );
  XNOR2_X1 U489 ( .A(n319), .B(b[5]), .ZN(n213) );
  OAI22_X1 U490 ( .A1(n293), .A2(n234), .B1(n336), .B2(n202), .ZN(n142) );
  XNOR2_X1 U491 ( .A(n310), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U492 ( .A(n319), .B(b[4]), .ZN(n214) );
  INV_X1 U493 ( .A(n336), .ZN(n143) );
  OAI22_X1 U494 ( .A1(n341), .A2(n209), .B1(n208), .B2(n336), .ZN(n174) );
  XNOR2_X1 U495 ( .A(n310), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U496 ( .A(n342), .B(n319), .ZN(n218) );
  XNOR2_X1 U497 ( .A(n310), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U498 ( .A(n310), .B(b[2]), .ZN(n216) );
  INV_X1 U499 ( .A(n319), .ZN(n243) );
  XNOR2_X1 U500 ( .A(n310), .B(b[1]), .ZN(n217) );
  XOR2_X1 U501 ( .A(n247), .B(n146), .Z(n231) );
  INV_X2 U502 ( .A(n146), .ZN(n255) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n35, n36, n38,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86, n87, n88,
         n91, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n139,
         n140, n142, n143, n145, n146, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n240, n241, n242, n243, n244, n245, n246, n247, n255, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n343, n344, n345, n346, n347, n348, n349, n350, n351;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n337), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n111), .B(n162), .CI(n156), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n164), .B(n170), .CI(n177), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n148), .B(n158), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n181), .B(n174), .CO(n134), .S(n135) );
  BUF_X1 U249 ( .A(n247), .Z(n328) );
  AND2_X1 U250 ( .A1(n99), .A2(n102), .ZN(n311) );
  BUF_X1 U251 ( .A(n247), .Z(n327) );
  INV_X1 U252 ( .A(n311), .ZN(n35) );
  AND3_X1 U253 ( .A1(n303), .A2(n304), .A3(n305), .ZN(product[15]) );
  OR2_X1 U254 ( .A1(n183), .A2(n151), .ZN(n286) );
  BUF_X2 U255 ( .A(n238), .Z(n346) );
  BUF_X1 U256 ( .A(n238), .Z(n345) );
  CLKBUF_X1 U257 ( .A(n55), .Z(n287) );
  INV_X1 U258 ( .A(n45), .ZN(n288) );
  CLKBUF_X1 U259 ( .A(n56), .Z(n289) );
  CLKBUF_X1 U260 ( .A(n350), .Z(n290) );
  OR2_X1 U261 ( .A1(n46), .A2(n41), .ZN(n291) );
  NOR2_X1 U262 ( .A1(n103), .A2(n106), .ZN(n292) );
  OAI21_X1 U263 ( .B1(n335), .B2(n16), .A(n17), .ZN(n15) );
  XNOR2_X1 U264 ( .A(n327), .B(n310), .ZN(n293) );
  CLKBUF_X1 U265 ( .A(n49), .Z(n294) );
  NOR2_X1 U266 ( .A1(n25), .A2(n20), .ZN(n295) );
  XNOR2_X1 U267 ( .A(n327), .B(a[2]), .ZN(n296) );
  CLKBUF_X1 U268 ( .A(n59), .Z(n297) );
  NOR2_X1 U269 ( .A1(n125), .A2(n128), .ZN(n59) );
  OAI21_X1 U270 ( .B1(n49), .B2(n291), .A(n38), .ZN(n298) );
  OAI21_X1 U271 ( .B1(n294), .B2(n291), .A(n38), .ZN(n299) );
  OAI21_X1 U272 ( .B1(n49), .B2(n291), .A(n38), .ZN(n36) );
  CLKBUF_X1 U273 ( .A(n73), .Z(n300) );
  CLKBUF_X1 U274 ( .A(n61), .Z(n301) );
  NOR2_X1 U275 ( .A1(n103), .A2(n106), .ZN(n41) );
  XOR2_X1 U276 ( .A(n152), .B(n94), .Z(n302) );
  XOR2_X1 U277 ( .A(n15), .B(n302), .Z(product[14]) );
  NAND2_X1 U278 ( .A1(n15), .A2(n152), .ZN(n303) );
  NAND2_X1 U279 ( .A1(n15), .A2(n94), .ZN(n304) );
  NAND2_X1 U280 ( .A1(n152), .A2(n94), .ZN(n305) );
  XNOR2_X1 U281 ( .A(n115), .B(n306), .ZN(n113) );
  XNOR2_X1 U282 ( .A(n117), .B(n120), .ZN(n306) );
  OR2_X1 U283 ( .A1(n133), .A2(n134), .ZN(n307) );
  NAND2_X1 U284 ( .A1(n293), .A2(n255), .ZN(n308) );
  NAND2_X1 U285 ( .A1(n293), .A2(n255), .ZN(n309) );
  NAND2_X1 U286 ( .A1(n231), .A2(n255), .ZN(n235) );
  INV_X1 U287 ( .A(n146), .ZN(n310) );
  AOI21_X1 U288 ( .B1(n341), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X1 U289 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  XNOR2_X1 U290 ( .A(n327), .B(n310), .ZN(n231) );
  INV_X2 U291 ( .A(n146), .ZN(n255) );
  OAI21_X1 U292 ( .B1(n52), .B2(n56), .A(n53), .ZN(n312) );
  XOR2_X1 U293 ( .A(n179), .B(n172), .Z(n313) );
  XOR2_X1 U294 ( .A(n131), .B(n313), .Z(n129) );
  NAND2_X1 U295 ( .A1(n131), .A2(n179), .ZN(n314) );
  NAND2_X1 U296 ( .A1(n131), .A2(n172), .ZN(n315) );
  NAND2_X1 U297 ( .A1(n179), .A2(n172), .ZN(n316) );
  NAND3_X1 U298 ( .A1(n314), .A2(n315), .A3(n316), .ZN(n128) );
  CLKBUF_X1 U299 ( .A(n246), .Z(n317) );
  NAND2_X1 U300 ( .A1(n115), .A2(n117), .ZN(n318) );
  NAND2_X1 U301 ( .A1(n115), .A2(n120), .ZN(n319) );
  NAND2_X1 U302 ( .A1(n117), .A2(n120), .ZN(n320) );
  NAND3_X1 U303 ( .A1(n318), .A2(n319), .A3(n320), .ZN(n112) );
  BUF_X2 U304 ( .A(n245), .Z(n321) );
  CLKBUF_X3 U305 ( .A(n236), .Z(n344) );
  NAND2_X1 U306 ( .A1(n246), .A2(n323), .ZN(n324) );
  NAND2_X1 U307 ( .A1(n322), .A2(a[2]), .ZN(n325) );
  NAND2_X1 U308 ( .A1(n324), .A2(n325), .ZN(n230) );
  INV_X1 U309 ( .A(n246), .ZN(n322) );
  INV_X1 U310 ( .A(a[2]), .ZN(n323) );
  OAI21_X1 U311 ( .B1(n292), .B2(n47), .A(n42), .ZN(n326) );
  NOR2_X1 U312 ( .A1(n113), .A2(n118), .ZN(n329) );
  XNOR2_X1 U313 ( .A(n246), .B(a[4]), .ZN(n330) );
  OAI21_X1 U314 ( .B1(n59), .B2(n61), .A(n60), .ZN(n331) );
  OAI21_X1 U315 ( .B1(n59), .B2(n61), .A(n60), .ZN(n332) );
  NAND2_X1 U316 ( .A1(n230), .A2(n296), .ZN(n333) );
  NAND2_X1 U317 ( .A1(n230), .A2(n296), .ZN(n334) );
  AOI21_X1 U318 ( .B1(n50), .B2(n331), .A(n51), .ZN(n335) );
  NAND2_X1 U319 ( .A1(n230), .A2(n296), .ZN(n234) );
  AOI21_X1 U320 ( .B1(n311), .B2(n338), .A(n28), .ZN(n336) );
  OAI22_X1 U321 ( .A1(n234), .A2(n203), .B1(n202), .B2(n346), .ZN(n337) );
  INV_X1 U322 ( .A(n326), .ZN(n38) );
  NAND2_X1 U323 ( .A1(n85), .A2(n288), .ZN(n5) );
  INV_X1 U324 ( .A(n46), .ZN(n85) );
  INV_X1 U325 ( .A(n47), .ZN(n45) );
  INV_X1 U326 ( .A(n65), .ZN(n63) );
  INV_X1 U327 ( .A(n77), .ZN(n75) );
  AOI21_X1 U328 ( .B1(n50), .B2(n332), .A(n312), .ZN(n49) );
  AOI21_X1 U329 ( .B1(n311), .B2(n338), .A(n28), .ZN(n26) );
  INV_X1 U330 ( .A(n30), .ZN(n28) );
  NOR2_X1 U331 ( .A1(n107), .A2(n112), .ZN(n46) );
  NAND2_X1 U332 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U333 ( .A(n297), .ZN(n88) );
  NAND2_X1 U334 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U335 ( .A(n20), .ZN(n81) );
  NAND2_X1 U336 ( .A1(n338), .A2(n30), .ZN(n2) );
  NAND2_X1 U337 ( .A1(n107), .A2(n112), .ZN(n47) );
  NOR2_X1 U338 ( .A1(n113), .A2(n118), .ZN(n52) );
  NAND2_X1 U339 ( .A1(n341), .A2(n65), .ZN(n9) );
  XOR2_X1 U340 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U341 ( .A1(n84), .A2(n42), .ZN(n4) );
  XNOR2_X1 U342 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U343 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U344 ( .B1(n57), .B2(n287), .A(n289), .ZN(n54) );
  INV_X1 U345 ( .A(n329), .ZN(n86) );
  NAND2_X1 U346 ( .A1(n113), .A2(n118), .ZN(n53) );
  XNOR2_X1 U347 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U348 ( .A1(n340), .A2(n77), .ZN(n12) );
  XOR2_X1 U349 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U350 ( .A1(n87), .A2(n289), .ZN(n7) );
  INV_X1 U351 ( .A(n287), .ZN(n87) );
  XNOR2_X1 U352 ( .A(n169), .B(n157), .ZN(n117) );
  OR2_X1 U353 ( .A1(n98), .A2(n97), .ZN(n338) );
  NOR2_X1 U354 ( .A1(n119), .A2(n124), .ZN(n55) );
  OR2_X1 U355 ( .A1(n169), .A2(n157), .ZN(n116) );
  NAND2_X1 U356 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U357 ( .A(n71), .ZN(n91) );
  INV_X1 U358 ( .A(n94), .ZN(n95) );
  NOR2_X1 U359 ( .A1(n96), .A2(n95), .ZN(n20) );
  XOR2_X1 U360 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U361 ( .A1(n307), .A2(n68), .ZN(n10) );
  NAND2_X1 U362 ( .A1(n119), .A2(n124), .ZN(n56) );
  OR2_X1 U363 ( .A1(n99), .A2(n102), .ZN(n339) );
  INV_X1 U364 ( .A(n80), .ZN(n78) );
  NAND2_X1 U365 ( .A1(n96), .A2(n95), .ZN(n21) );
  OR2_X1 U366 ( .A1(n182), .A2(n175), .ZN(n340) );
  OR2_X1 U367 ( .A1(n129), .A2(n132), .ZN(n341) );
  NAND2_X1 U368 ( .A1(n125), .A2(n128), .ZN(n60) );
  AND2_X1 U369 ( .A1(n351), .A2(n143), .ZN(n175) );
  AND2_X1 U370 ( .A1(n351), .A2(n140), .ZN(n167) );
  OR2_X1 U371 ( .A1(n351), .A2(n241), .ZN(n201) );
  BUF_X1 U372 ( .A(n227), .Z(n351) );
  INV_X1 U373 ( .A(n139), .ZN(n160) );
  AND2_X1 U374 ( .A1(n351), .A2(n137), .ZN(n159) );
  NOR2_X1 U375 ( .A1(n133), .A2(n134), .ZN(n67) );
  INV_X1 U376 ( .A(n100), .ZN(n101) );
  INV_X1 U377 ( .A(n142), .ZN(n168) );
  INV_X1 U378 ( .A(n136), .ZN(n152) );
  NAND2_X1 U379 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U380 ( .A1(n351), .A2(n240), .ZN(n192) );
  AND2_X1 U381 ( .A1(n286), .A2(n80), .ZN(product[1]) );
  OR2_X1 U382 ( .A1(n351), .A2(n243), .ZN(n219) );
  OR2_X1 U383 ( .A1(n351), .A2(n242), .ZN(n210) );
  AND2_X1 U384 ( .A1(n351), .A2(n146), .ZN(product[0]) );
  OAI21_X1 U385 ( .B1(n297), .B2(n301), .A(n60), .ZN(n58) );
  NAND2_X1 U386 ( .A1(n182), .A2(n175), .ZN(n77) );
  CLKBUF_X1 U387 ( .A(n236), .Z(n343) );
  XNOR2_X1 U388 ( .A(n245), .B(a[6]), .ZN(n236) );
  XNOR2_X1 U389 ( .A(n327), .B(a[2]), .ZN(n238) );
  XNOR2_X1 U390 ( .A(n246), .B(a[4]), .ZN(n237) );
  INV_X1 U391 ( .A(n70), .ZN(n69) );
  INV_X1 U392 ( .A(n244), .ZN(n240) );
  XNOR2_X1 U393 ( .A(n351), .B(n244), .ZN(n191) );
  XNOR2_X1 U394 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U395 ( .A(n244), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U396 ( .A(n244), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U397 ( .A(n244), .B(b[5]), .ZN(n186) );
  XOR2_X1 U398 ( .A(n244), .B(a[6]), .Z(n228) );
  NAND2_X1 U399 ( .A1(n183), .A2(n151), .ZN(n80) );
  OAI22_X1 U400 ( .A1(n309), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U401 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U402 ( .A1(n308), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U403 ( .A1(n309), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  OAI22_X1 U404 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OAI22_X1 U405 ( .A1(n309), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OAI22_X1 U406 ( .A1(n308), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U407 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  NOR2_X1 U408 ( .A1(n25), .A2(n20), .ZN(n18) );
  INV_X1 U409 ( .A(n25), .ZN(n23) );
  NAND2_X1 U410 ( .A1(n229), .A2(n330), .ZN(n347) );
  NAND2_X1 U411 ( .A1(n229), .A2(n330), .ZN(n348) );
  CLKBUF_X1 U412 ( .A(n237), .Z(n349) );
  NAND2_X1 U413 ( .A1(n229), .A2(n237), .ZN(n233) );
  INV_X1 U414 ( .A(n292), .ZN(n84) );
  NOR2_X1 U415 ( .A1(n46), .A2(n41), .ZN(n39) );
  OAI21_X1 U416 ( .B1(n41), .B2(n47), .A(n42), .ZN(n40) );
  NAND2_X1 U417 ( .A1(n103), .A2(n106), .ZN(n42) );
  INV_X1 U418 ( .A(n110), .ZN(n111) );
  NAND2_X1 U419 ( .A1(n129), .A2(n132), .ZN(n65) );
  XNOR2_X1 U420 ( .A(n244), .B(b[6]), .ZN(n185) );
  INV_X1 U421 ( .A(n145), .ZN(n176) );
  OAI22_X1 U422 ( .A1(n211), .A2(n308), .B1(n211), .B2(n255), .ZN(n145) );
  NAND2_X1 U423 ( .A1(n228), .A2(n344), .ZN(n350) );
  NAND2_X1 U424 ( .A1(n228), .A2(n343), .ZN(n232) );
  XOR2_X1 U425 ( .A(n245), .B(a[4]), .Z(n229) );
  INV_X1 U426 ( .A(n245), .ZN(n241) );
  XNOR2_X1 U427 ( .A(n321), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U428 ( .A(n321), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U429 ( .A(n321), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U430 ( .A(n321), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U431 ( .A(n321), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U432 ( .A(n351), .B(n321), .ZN(n200) );
  XNOR2_X1 U433 ( .A(n9), .B(n66), .ZN(product[5]) );
  OAI21_X1 U434 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  XOR2_X1 U435 ( .A(n11), .B(n300), .Z(product[3]) );
  AOI21_X1 U436 ( .B1(n340), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U437 ( .A(n336), .ZN(n24) );
  OAI21_X1 U438 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  NAND2_X1 U439 ( .A1(n98), .A2(n97), .ZN(n30) );
  XNOR2_X1 U440 ( .A(n244), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U441 ( .A(n321), .B(b[7]), .ZN(n193) );
  OAI22_X1 U442 ( .A1(n184), .A2(n290), .B1(n184), .B2(n344), .ZN(n136) );
  OAI22_X1 U443 ( .A1(n290), .A2(n185), .B1(n184), .B2(n344), .ZN(n94) );
  OAI22_X1 U444 ( .A1(n290), .A2(n188), .B1(n187), .B2(n344), .ZN(n155) );
  OAI22_X1 U445 ( .A1(n290), .A2(n187), .B1(n186), .B2(n344), .ZN(n154) );
  OAI22_X1 U446 ( .A1(n350), .A2(n190), .B1(n189), .B2(n344), .ZN(n157) );
  OAI22_X1 U447 ( .A1(n350), .A2(n186), .B1(n185), .B2(n344), .ZN(n153) );
  INV_X1 U448 ( .A(n344), .ZN(n137) );
  OAI22_X1 U449 ( .A1(n350), .A2(n189), .B1(n188), .B2(n344), .ZN(n156) );
  OAI22_X1 U450 ( .A1(n232), .A2(n240), .B1(n192), .B2(n344), .ZN(n148) );
  OAI22_X1 U451 ( .A1(n232), .A2(n191), .B1(n190), .B2(n344), .ZN(n158) );
  NAND2_X1 U452 ( .A1(n339), .A2(n338), .ZN(n25) );
  NAND2_X1 U453 ( .A1(n339), .A2(n35), .ZN(n3) );
  OAI21_X1 U454 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  NOR2_X1 U455 ( .A1(n329), .A2(n55), .ZN(n50) );
  NAND2_X1 U456 ( .A1(n39), .A2(n18), .ZN(n16) );
  AOI21_X1 U457 ( .B1(n40), .B2(n295), .A(n19), .ZN(n17) );
  XOR2_X1 U458 ( .A(n22), .B(n1), .Z(product[13]) );
  INV_X1 U459 ( .A(n58), .ZN(n57) );
  OAI22_X1 U460 ( .A1(n347), .A2(n199), .B1(n198), .B2(n349), .ZN(n165) );
  OAI22_X1 U461 ( .A1(n347), .A2(n197), .B1(n196), .B2(n237), .ZN(n163) );
  OAI22_X1 U462 ( .A1(n348), .A2(n198), .B1(n197), .B2(n237), .ZN(n164) );
  OAI22_X1 U463 ( .A1(n348), .A2(n194), .B1(n193), .B2(n349), .ZN(n100) );
  OAI22_X1 U464 ( .A1(n348), .A2(n196), .B1(n195), .B2(n237), .ZN(n162) );
  INV_X1 U465 ( .A(n330), .ZN(n140) );
  OAI22_X1 U466 ( .A1(n193), .A2(n347), .B1(n193), .B2(n349), .ZN(n139) );
  OAI22_X1 U467 ( .A1(n233), .A2(n241), .B1(n201), .B2(n237), .ZN(n149) );
  OAI22_X1 U468 ( .A1(n347), .A2(n195), .B1(n194), .B2(n330), .ZN(n161) );
  OAI22_X1 U469 ( .A1(n233), .A2(n200), .B1(n199), .B2(n237), .ZN(n166) );
  INV_X1 U470 ( .A(n317), .ZN(n242) );
  XNOR2_X1 U471 ( .A(n246), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U472 ( .A(n246), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U473 ( .A(n246), .B(b[5]), .ZN(n204) );
  XNOR2_X1 U474 ( .A(n351), .B(n317), .ZN(n209) );
  XNOR2_X1 U475 ( .A(n246), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U476 ( .A(n246), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U477 ( .A(n246), .B(b[7]), .ZN(n202) );
  XOR2_X1 U478 ( .A(n31), .B(n2), .Z(product[12]) );
  XNOR2_X1 U479 ( .A(n328), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U480 ( .A(n328), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U481 ( .A(n328), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U482 ( .A(n328), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U483 ( .A(n328), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U484 ( .A(n351), .B(n328), .ZN(n218) );
  XNOR2_X1 U485 ( .A(n328), .B(b[1]), .ZN(n217) );
  INV_X1 U486 ( .A(n328), .ZN(n243) );
  XNOR2_X1 U487 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U488 ( .A(n8), .B(n301), .Z(product[6]) );
  AOI21_X1 U489 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  NOR2_X1 U490 ( .A1(n135), .A2(n150), .ZN(n71) );
  NAND2_X1 U491 ( .A1(n135), .A2(n150), .ZN(n72) );
  XNOR2_X1 U492 ( .A(n317), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U493 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U494 ( .A(n321), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U495 ( .A(n328), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U496 ( .A(n299), .B(n3), .ZN(product[11]) );
  AOI21_X1 U497 ( .B1(n298), .B2(n339), .A(n311), .ZN(n31) );
  AOI21_X1 U498 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U499 ( .A(n335), .ZN(n48) );
  OAI22_X1 U500 ( .A1(n333), .A2(n204), .B1(n203), .B2(n346), .ZN(n169) );
  OAI22_X1 U501 ( .A1(n334), .A2(n207), .B1(n206), .B2(n345), .ZN(n172) );
  OAI22_X1 U502 ( .A1(n333), .A2(n206), .B1(n205), .B2(n346), .ZN(n171) );
  OAI22_X1 U503 ( .A1(n334), .A2(n205), .B1(n204), .B2(n345), .ZN(n170) );
  OAI22_X1 U504 ( .A1(n334), .A2(n208), .B1(n207), .B2(n346), .ZN(n173) );
  OAI22_X1 U505 ( .A1(n333), .A2(n242), .B1(n210), .B2(n345), .ZN(n150) );
  OAI22_X1 U506 ( .A1(n333), .A2(n203), .B1(n202), .B2(n346), .ZN(n110) );
  OAI22_X1 U507 ( .A1(n202), .A2(n234), .B1(n202), .B2(n346), .ZN(n142) );
  INV_X1 U508 ( .A(n346), .ZN(n143) );
  OAI22_X1 U509 ( .A1(n234), .A2(n209), .B1(n208), .B2(n345), .ZN(n174) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n75, n77, n78, n80, n81, n84, n85, n86,
         n87, n88, n90, n91, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n142, n143, n145, n146, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n227, n228, n229, n232, n233, n234, n235, n236,
         n237, n238, n240, n241, n242, n243, n244, n245, n246, n247, n255,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n161), .B(n110), .CI(n168), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n162), .B(n156), .CI(n111), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n177), .B(n170), .CI(n164), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n149), .B(n166), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  OR2_X1 U249 ( .A1(n98), .A2(n97), .ZN(n285) );
  OR2_X1 U250 ( .A1(n183), .A2(n151), .ZN(n286) );
  INV_X1 U251 ( .A(n240), .ZN(n287) );
  XNOR2_X1 U252 ( .A(n115), .B(n303), .ZN(n288) );
  OAI21_X2 U253 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  XNOR2_X1 U254 ( .A(n292), .B(b[4]), .ZN(n289) );
  BUF_X2 U255 ( .A(n238), .Z(n290) );
  CLKBUF_X1 U256 ( .A(n238), .Z(n337) );
  AOI21_X2 U257 ( .B1(n336), .B2(n66), .A(n63), .ZN(n291) );
  AOI21_X1 U258 ( .B1(n336), .B2(n66), .A(n63), .ZN(n61) );
  BUF_X2 U259 ( .A(n246), .Z(n292) );
  CLKBUF_X1 U260 ( .A(n234), .Z(n293) );
  OAI21_X1 U261 ( .B1(n59), .B2(n291), .A(n60), .ZN(n294) );
  AOI21_X1 U262 ( .B1(n320), .B2(n285), .A(n28), .ZN(n295) );
  CLKBUF_X1 U263 ( .A(n291), .Z(n296) );
  CLKBUF_X1 U264 ( .A(n55), .Z(n297) );
  NOR2_X1 U265 ( .A1(n103), .A2(n106), .ZN(n298) );
  AND2_X1 U266 ( .A1(n102), .A2(n99), .ZN(n320) );
  CLKBUF_X1 U267 ( .A(n245), .Z(n304) );
  BUF_X2 U268 ( .A(n245), .Z(n317) );
  OR2_X2 U269 ( .A1(n299), .A2(n146), .ZN(n235) );
  XNOR2_X1 U270 ( .A(n247), .B(n146), .ZN(n299) );
  OAI21_X1 U271 ( .B1(n59), .B2(n291), .A(n60), .ZN(n300) );
  CLKBUF_X1 U272 ( .A(n178), .Z(n301) );
  INV_X1 U273 ( .A(n146), .ZN(n255) );
  CLKBUF_X1 U274 ( .A(n56), .Z(n302) );
  INV_X1 U275 ( .A(n320), .ZN(n35) );
  XNOR2_X1 U276 ( .A(n115), .B(n303), .ZN(n113) );
  XNOR2_X1 U277 ( .A(n120), .B(n117), .ZN(n303) );
  BUF_X2 U278 ( .A(n237), .Z(n338) );
  OAI21_X1 U279 ( .B1(n330), .B2(n37), .A(n38), .ZN(n36) );
  NAND2_X1 U280 ( .A1(n237), .A2(n229), .ZN(n305) );
  NAND2_X1 U281 ( .A1(n237), .A2(n229), .ZN(n233) );
  BUF_X1 U282 ( .A(n236), .Z(n343) );
  BUF_X2 U283 ( .A(n247), .Z(n306) );
  INV_X1 U284 ( .A(n323), .ZN(n307) );
  CLKBUF_X1 U285 ( .A(n237), .Z(n339) );
  NAND2_X1 U286 ( .A1(n115), .A2(n120), .ZN(n308) );
  NAND2_X1 U287 ( .A1(n115), .A2(n117), .ZN(n309) );
  NAND2_X1 U288 ( .A1(n120), .A2(n117), .ZN(n310) );
  NAND3_X1 U289 ( .A1(n308), .A2(n309), .A3(n310), .ZN(n112) );
  NAND2_X1 U290 ( .A1(n238), .A2(n332), .ZN(n311) );
  OAI22_X1 U291 ( .A1(n293), .A2(n206), .B1(n289), .B2(n290), .ZN(n312) );
  NAND2_X1 U292 ( .A1(n238), .A2(n332), .ZN(n234) );
  XOR2_X1 U293 ( .A(n171), .B(n178), .Z(n313) );
  XOR2_X1 U294 ( .A(n159), .B(n313), .Z(n127) );
  NAND2_X1 U295 ( .A1(n159), .A2(n301), .ZN(n314) );
  NAND2_X1 U296 ( .A1(n159), .A2(n312), .ZN(n315) );
  NAND2_X1 U297 ( .A1(n301), .A2(n312), .ZN(n316) );
  NAND3_X1 U298 ( .A1(n314), .A2(n315), .A3(n316), .ZN(n126) );
  OAI21_X1 U299 ( .B1(n41), .B2(n47), .A(n42), .ZN(n318) );
  CLKBUF_X1 U300 ( .A(n340), .Z(n319) );
  CLKBUF_X1 U301 ( .A(n247), .Z(n321) );
  NOR2_X1 U302 ( .A1(n113), .A2(n118), .ZN(n322) );
  NOR2_X1 U303 ( .A1(n288), .A2(n118), .ZN(n52) );
  NOR2_X2 U304 ( .A1(n125), .A2(n128), .ZN(n59) );
  NAND2_X1 U305 ( .A1(n246), .A2(n324), .ZN(n325) );
  NAND2_X1 U306 ( .A1(n323), .A2(a[2]), .ZN(n326) );
  NAND2_X1 U307 ( .A1(n325), .A2(n326), .ZN(n332) );
  INV_X1 U308 ( .A(n246), .ZN(n323) );
  INV_X1 U309 ( .A(a[2]), .ZN(n324) );
  OAI21_X1 U310 ( .B1(n322), .B2(n56), .A(n53), .ZN(n327) );
  CLKBUF_X1 U311 ( .A(n36), .Z(n328) );
  BUF_X1 U312 ( .A(n236), .Z(n341) );
  OAI21_X1 U313 ( .B1(n59), .B2(n296), .A(n60), .ZN(n329) );
  AOI21_X1 U314 ( .B1(n300), .B2(n50), .A(n51), .ZN(n330) );
  AOI21_X1 U315 ( .B1(n58), .B2(n50), .A(n327), .ZN(n331) );
  NOR2_X1 U316 ( .A1(n119), .A2(n124), .ZN(n55) );
  NAND2_X1 U317 ( .A1(n119), .A2(n124), .ZN(n56) );
  INV_X1 U318 ( .A(n39), .ZN(n37) );
  INV_X1 U319 ( .A(n318), .ZN(n38) );
  NAND2_X1 U320 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U321 ( .A(n295), .ZN(n24) );
  INV_X1 U322 ( .A(n25), .ZN(n23) );
  INV_X1 U323 ( .A(n47), .ZN(n45) );
  AOI21_X1 U324 ( .B1(n320), .B2(n285), .A(n28), .ZN(n26) );
  INV_X1 U325 ( .A(n30), .ZN(n28) );
  AOI21_X1 U326 ( .B1(n333), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U327 ( .A(n77), .ZN(n75) );
  NAND2_X1 U328 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U329 ( .A(n59), .ZN(n88) );
  NAND2_X1 U330 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U331 ( .A(n20), .ZN(n81) );
  NAND2_X1 U332 ( .A1(n285), .A2(n30), .ZN(n2) );
  XOR2_X1 U333 ( .A(n43), .B(n4), .Z(product[10]) );
  NAND2_X1 U334 ( .A1(n84), .A2(n42), .ZN(n4) );
  INV_X1 U335 ( .A(n298), .ZN(n84) );
  INV_X1 U336 ( .A(n80), .ZN(n78) );
  XNOR2_X1 U337 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U338 ( .A1(n86), .A2(n53), .ZN(n6) );
  OAI21_X1 U339 ( .B1(n57), .B2(n297), .A(n302), .ZN(n54) );
  XNOR2_X1 U340 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U341 ( .A1(n333), .A2(n77), .ZN(n12) );
  NAND2_X1 U342 ( .A1(n107), .A2(n112), .ZN(n47) );
  XOR2_X1 U343 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U344 ( .A1(n87), .A2(n302), .ZN(n7) );
  INV_X1 U345 ( .A(n297), .ZN(n87) );
  NOR2_X1 U346 ( .A1(n103), .A2(n106), .ZN(n41) );
  OR2_X1 U347 ( .A1(n169), .A2(n157), .ZN(n116) );
  NAND2_X1 U348 ( .A1(n91), .A2(n72), .ZN(n11) );
  INV_X1 U349 ( .A(n71), .ZN(n91) );
  XNOR2_X1 U350 ( .A(n169), .B(n157), .ZN(n117) );
  INV_X1 U351 ( .A(n94), .ZN(n95) );
  NOR2_X1 U352 ( .A1(n96), .A2(n95), .ZN(n20) );
  XOR2_X1 U353 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U354 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U355 ( .A(n67), .ZN(n90) );
  INV_X1 U356 ( .A(n70), .ZN(n69) );
  OR2_X1 U357 ( .A1(n182), .A2(n175), .ZN(n333) );
  NAND2_X1 U358 ( .A1(n125), .A2(n128), .ZN(n60) );
  NAND2_X1 U359 ( .A1(n96), .A2(n95), .ZN(n21) );
  NAND2_X1 U360 ( .A1(n103), .A2(n106), .ZN(n42) );
  AND2_X1 U361 ( .A1(n286), .A2(n80), .ZN(product[1]) );
  OR2_X1 U362 ( .A1(n99), .A2(n102), .ZN(n335) );
  AND2_X1 U363 ( .A1(n344), .A2(n143), .ZN(n175) );
  OR2_X1 U364 ( .A1(n129), .A2(n132), .ZN(n336) );
  INV_X1 U365 ( .A(n14), .ZN(product[15]) );
  AND2_X1 U366 ( .A1(n344), .A2(n140), .ZN(n167) );
  OAI22_X1 U367 ( .A1(n235), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U368 ( .A1(n235), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  OAI22_X1 U369 ( .A1(n235), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  OAI22_X1 U370 ( .A1(n235), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OR2_X1 U371 ( .A1(n344), .A2(n243), .ZN(n219) );
  OR2_X1 U372 ( .A1(n344), .A2(n241), .ZN(n201) );
  NOR2_X1 U373 ( .A1(n133), .A2(n134), .ZN(n67) );
  BUF_X1 U374 ( .A(n227), .Z(n344) );
  INV_X1 U375 ( .A(n139), .ZN(n160) );
  OAI22_X1 U376 ( .A1(n235), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  AND2_X1 U377 ( .A1(n344), .A2(n137), .ZN(n159) );
  OAI22_X1 U378 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  INV_X1 U379 ( .A(n100), .ZN(n101) );
  INV_X1 U380 ( .A(n136), .ZN(n152) );
  NAND2_X1 U381 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U382 ( .A1(n344), .A2(n240), .ZN(n192) );
  OR2_X1 U383 ( .A1(n344), .A2(n242), .ZN(n210) );
  OAI22_X1 U384 ( .A1(n235), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  XNOR2_X1 U385 ( .A(n287), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U386 ( .A(n244), .B(b[6]), .ZN(n185) );
  XNOR2_X1 U387 ( .A(n287), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U388 ( .A(n244), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U389 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U390 ( .A(n344), .B(n244), .ZN(n191) );
  INV_X1 U391 ( .A(n244), .ZN(n240) );
  AND2_X1 U392 ( .A1(n344), .A2(n146), .ZN(product[0]) );
  XNOR2_X1 U393 ( .A(n247), .B(a[2]), .ZN(n238) );
  XNOR2_X1 U394 ( .A(n246), .B(a[4]), .ZN(n237) );
  NAND2_X1 U395 ( .A1(n335), .A2(n35), .ZN(n3) );
  OAI21_X1 U396 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  NAND2_X1 U397 ( .A1(n228), .A2(n341), .ZN(n340) );
  BUF_X2 U398 ( .A(n341), .Z(n342) );
  NAND2_X1 U399 ( .A1(n228), .A2(n236), .ZN(n232) );
  XNOR2_X1 U400 ( .A(n245), .B(a[6]), .ZN(n236) );
  INV_X1 U401 ( .A(n110), .ZN(n111) );
  NAND2_X1 U402 ( .A1(n98), .A2(n97), .ZN(n30) );
  INV_X1 U403 ( .A(n46), .ZN(n85) );
  NOR2_X1 U404 ( .A1(n46), .A2(n41), .ZN(n39) );
  NOR2_X1 U405 ( .A1(n107), .A2(n112), .ZN(n46) );
  NAND2_X1 U406 ( .A1(n288), .A2(n118), .ZN(n53) );
  XNOR2_X1 U407 ( .A(n9), .B(n66), .ZN(product[5]) );
  NAND2_X1 U408 ( .A1(n182), .A2(n175), .ZN(n77) );
  INV_X1 U409 ( .A(n65), .ZN(n63) );
  NAND2_X1 U410 ( .A1(n336), .A2(n65), .ZN(n9) );
  OAI21_X1 U411 ( .B1(n298), .B2(n47), .A(n42), .ZN(n40) );
  INV_X1 U412 ( .A(n145), .ZN(n176) );
  OAI22_X1 U413 ( .A1(n211), .A2(n235), .B1(n211), .B2(n255), .ZN(n145) );
  OAI22_X1 U414 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  XOR2_X1 U415 ( .A(n244), .B(a[6]), .Z(n228) );
  NAND2_X1 U416 ( .A1(n129), .A2(n132), .ZN(n65) );
  NOR2_X1 U417 ( .A1(n135), .A2(n150), .ZN(n71) );
  OAI22_X1 U418 ( .A1(n184), .A2(n319), .B1(n184), .B2(n342), .ZN(n136) );
  OAI22_X1 U419 ( .A1(n319), .A2(n185), .B1(n184), .B2(n343), .ZN(n94) );
  OAI22_X1 U420 ( .A1(n319), .A2(n188), .B1(n187), .B2(n342), .ZN(n155) );
  OAI22_X1 U421 ( .A1(n340), .A2(n187), .B1(n186), .B2(n343), .ZN(n154) );
  OAI22_X1 U422 ( .A1(n340), .A2(n186), .B1(n185), .B2(n342), .ZN(n153) );
  OAI22_X1 U423 ( .A1(n340), .A2(n190), .B1(n189), .B2(n343), .ZN(n157) );
  OAI22_X1 U424 ( .A1(n340), .A2(n189), .B1(n188), .B2(n342), .ZN(n156) );
  INV_X1 U425 ( .A(n342), .ZN(n137) );
  OAI22_X1 U426 ( .A1(n232), .A2(n240), .B1(n192), .B2(n343), .ZN(n148) );
  OAI22_X1 U427 ( .A1(n232), .A2(n191), .B1(n190), .B2(n343), .ZN(n158) );
  XNOR2_X1 U428 ( .A(b[3]), .B(n317), .ZN(n197) );
  XNOR2_X1 U429 ( .A(n317), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U430 ( .A(n317), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U431 ( .A(n317), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U432 ( .A(n304), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U433 ( .A(n344), .B(n317), .ZN(n200) );
  INV_X1 U434 ( .A(n304), .ZN(n241) );
  XOR2_X1 U435 ( .A(n245), .B(a[4]), .Z(n229) );
  XNOR2_X1 U436 ( .A(n317), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U437 ( .A(n244), .B(b[2]), .ZN(n189) );
  OAI21_X1 U438 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  INV_X1 U439 ( .A(n142), .ZN(n168) );
  XOR2_X1 U440 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U441 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  NAND2_X1 U442 ( .A1(n183), .A2(n151), .ZN(n80) );
  AOI21_X1 U443 ( .B1(n294), .B2(n50), .A(n327), .ZN(n49) );
  AOI21_X1 U444 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  INV_X1 U445 ( .A(n52), .ZN(n86) );
  NOR2_X1 U446 ( .A1(n52), .A2(n55), .ZN(n50) );
  OAI21_X1 U447 ( .B1(n322), .B2(n56), .A(n53), .ZN(n51) );
  XOR2_X1 U448 ( .A(n22), .B(n1), .Z(product[13]) );
  NOR2_X1 U449 ( .A1(n25), .A2(n20), .ZN(n18) );
  NAND2_X1 U450 ( .A1(n335), .A2(n285), .ZN(n25) );
  NAND2_X1 U451 ( .A1(n39), .A2(n18), .ZN(n16) );
  XOR2_X1 U452 ( .A(n31), .B(n2), .Z(product[12]) );
  INV_X1 U453 ( .A(n329), .ZN(n57) );
  NAND2_X1 U454 ( .A1(n135), .A2(n150), .ZN(n72) );
  XNOR2_X1 U455 ( .A(n48), .B(n5), .ZN(product[9]) );
  XOR2_X1 U456 ( .A(n8), .B(n296), .Z(product[6]) );
  AOI21_X1 U457 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  OAI22_X1 U458 ( .A1(n305), .A2(n199), .B1(n198), .B2(n338), .ZN(n165) );
  OAI22_X1 U459 ( .A1(n305), .A2(n197), .B1(n196), .B2(n339), .ZN(n163) );
  OAI22_X1 U460 ( .A1(n305), .A2(n194), .B1(n193), .B2(n339), .ZN(n100) );
  OAI22_X1 U461 ( .A1(n305), .A2(n196), .B1(n195), .B2(n338), .ZN(n162) );
  OAI22_X1 U462 ( .A1(n305), .A2(n198), .B1(n197), .B2(n339), .ZN(n164) );
  OAI22_X1 U463 ( .A1(n193), .A2(n305), .B1(n193), .B2(n338), .ZN(n139) );
  OAI22_X1 U464 ( .A1(n233), .A2(n195), .B1(n194), .B2(n338), .ZN(n161) );
  INV_X1 U465 ( .A(n339), .ZN(n140) );
  OAI22_X1 U466 ( .A1(n233), .A2(n241), .B1(n201), .B2(n338), .ZN(n149) );
  XNOR2_X1 U467 ( .A(n292), .B(b[3]), .ZN(n206) );
  OAI22_X1 U468 ( .A1(n233), .A2(n200), .B1(n199), .B2(n338), .ZN(n166) );
  XNOR2_X1 U469 ( .A(n292), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U470 ( .A(n307), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U471 ( .A(n307), .B(b[5]), .ZN(n204) );
  INV_X1 U472 ( .A(n307), .ZN(n242) );
  XNOR2_X1 U473 ( .A(n292), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U474 ( .A(n292), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U475 ( .A(n344), .B(n307), .ZN(n209) );
  XNOR2_X1 U476 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U477 ( .A(n304), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U478 ( .A(n307), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U479 ( .A(n328), .B(n3), .ZN(product[11]) );
  AOI21_X1 U480 ( .B1(n36), .B2(n335), .A(n320), .ZN(n31) );
  AOI21_X1 U481 ( .B1(n36), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U482 ( .B1(n331), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U483 ( .A(n49), .ZN(n48) );
  OAI22_X1 U484 ( .A1(n311), .A2(n204), .B1(n203), .B2(n290), .ZN(n169) );
  OAI22_X1 U485 ( .A1(n311), .A2(n207), .B1(n206), .B2(n290), .ZN(n172) );
  OAI22_X1 U486 ( .A1(n206), .A2(n234), .B1(n205), .B2(n337), .ZN(n171) );
  OAI22_X1 U487 ( .A1(n311), .A2(n289), .B1(n204), .B2(n290), .ZN(n170) );
  OAI22_X1 U488 ( .A1(n311), .A2(n208), .B1(n207), .B2(n290), .ZN(n173) );
  OAI22_X1 U489 ( .A1(n311), .A2(n242), .B1(n210), .B2(n290), .ZN(n150) );
  OAI22_X1 U490 ( .A1(n234), .A2(n203), .B1(n202), .B2(n337), .ZN(n110) );
  XNOR2_X1 U491 ( .A(n306), .B(b[5]), .ZN(n213) );
  OAI22_X1 U492 ( .A1(n202), .A2(n234), .B1(n202), .B2(n337), .ZN(n142) );
  XNOR2_X1 U493 ( .A(n321), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U494 ( .A(n306), .B(b[4]), .ZN(n214) );
  INV_X1 U495 ( .A(n290), .ZN(n143) );
  OAI22_X1 U496 ( .A1(n311), .A2(n209), .B1(n208), .B2(n290), .ZN(n174) );
  XNOR2_X1 U497 ( .A(n321), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U498 ( .A(n344), .B(n321), .ZN(n218) );
  XNOR2_X1 U499 ( .A(n321), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U500 ( .A(n306), .B(b[2]), .ZN(n216) );
  INV_X1 U501 ( .A(n306), .ZN(n243) );
  XNOR2_X1 U502 ( .A(n306), .B(b[1]), .ZN(n217) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1_DW_mult_tc_1 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n24, n25, n26, n30, n31, n35, n36, n38, n39,
         n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n75, n77, n78, n80, n81, n85, n87, n88, n90, n91, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n139, n140,
         n142, n143, n145, n146, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n240, n241, n242, n243, n244, n245, n246, n247, n255, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n340, n341, n342,
         n343, n344, n345, n346, n347;
  assign n146 = a[0];
  assign n227 = b[0];
  assign n244 = a[7];
  assign n245 = a[5];
  assign n246 = a[3];
  assign n247 = a[1];

  FA_X1 U2 ( .A(n152), .B(n94), .CI(n15), .CO(n14), .S(product[14]) );
  FA_X1 U109 ( .A(n153), .B(n100), .CI(n160), .CO(n96), .S(n97) );
  FA_X1 U110 ( .A(n101), .B(n154), .CI(n104), .CO(n98), .S(n99) );
  FA_X1 U112 ( .A(n108), .B(n155), .CI(n105), .CO(n102), .S(n103) );
  FA_X1 U113 ( .A(n168), .B(n329), .CI(n161), .CO(n104), .S(n105) );
  FA_X1 U114 ( .A(n114), .B(n116), .CI(n109), .CO(n106), .S(n107) );
  FA_X1 U115 ( .A(n162), .B(n111), .CI(n156), .CO(n108), .S(n109) );
  FA_X1 U118 ( .A(n176), .B(n163), .CI(n122), .CO(n114), .S(n115) );
  FA_X1 U121 ( .A(n126), .B(n123), .CI(n121), .CO(n118), .S(n119) );
  FA_X1 U122 ( .A(n164), .B(n177), .CI(n170), .CO(n120), .S(n121) );
  HA_X1 U123 ( .A(n158), .B(n148), .CO(n122), .S(n123) );
  FA_X1 U124 ( .A(n130), .B(n165), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U125 ( .A(n178), .B(n159), .CI(n171), .CO(n126), .S(n127) );
  FA_X1 U126 ( .A(n172), .B(n179), .CI(n131), .CO(n128), .S(n129) );
  HA_X1 U127 ( .A(n166), .B(n149), .CO(n130), .S(n131) );
  FA_X1 U128 ( .A(n180), .B(n167), .CI(n173), .CO(n132), .S(n133) );
  HA_X1 U129 ( .A(n174), .B(n181), .CO(n134), .S(n135) );
  CLKBUF_X3 U249 ( .A(n246), .Z(n312) );
  BUF_X1 U250 ( .A(n236), .Z(n343) );
  CLKBUF_X2 U251 ( .A(n247), .Z(n309) );
  OAI21_X1 U252 ( .B1(n52), .B2(n56), .A(n53), .ZN(n285) );
  NAND2_X1 U253 ( .A1(n303), .A2(n307), .ZN(n334) );
  INV_X1 U254 ( .A(n293), .ZN(n30) );
  OR2_X1 U255 ( .A1(n103), .A2(n106), .ZN(n286) );
  OR2_X1 U256 ( .A1(n183), .A2(n151), .ZN(n287) );
  AND2_X1 U257 ( .A1(n98), .A2(n97), .ZN(n293) );
  OR2_X1 U258 ( .A1(n46), .A2(n41), .ZN(n288) );
  CLKBUF_X1 U259 ( .A(n245), .Z(n289) );
  XNOR2_X1 U260 ( .A(n309), .B(b[7]), .ZN(n290) );
  CLKBUF_X1 U261 ( .A(n245), .Z(n291) );
  NAND2_X1 U262 ( .A1(n231), .A2(n255), .ZN(n292) );
  NAND2_X1 U263 ( .A1(n231), .A2(n255), .ZN(n235) );
  XNOR2_X1 U264 ( .A(n169), .B(n157), .ZN(n117) );
  OAI21_X1 U265 ( .B1(n59), .B2(n61), .A(n60), .ZN(n294) );
  INV_X1 U266 ( .A(n35), .ZN(n295) );
  INV_X1 U267 ( .A(n315), .ZN(n35) );
  AND2_X1 U268 ( .A1(n102), .A2(n99), .ZN(n315) );
  AND2_X1 U269 ( .A1(n337), .A2(n336), .ZN(n296) );
  OR2_X2 U270 ( .A1(n98), .A2(n97), .ZN(n336) );
  BUF_X1 U271 ( .A(n327), .Z(n297) );
  BUF_X1 U272 ( .A(n327), .Z(n298) );
  XNOR2_X1 U273 ( .A(n246), .B(a[4]), .ZN(n327) );
  CLKBUF_X1 U274 ( .A(n341), .Z(n299) );
  CLKBUF_X1 U275 ( .A(n245), .Z(n300) );
  NOR2_X1 U276 ( .A1(n103), .A2(n106), .ZN(n301) );
  NOR2_X1 U277 ( .A1(n103), .A2(n106), .ZN(n41) );
  NOR2_X1 U278 ( .A1(n25), .A2(n20), .ZN(n302) );
  XOR2_X1 U279 ( .A(n244), .B(a[6]), .Z(n303) );
  CLKBUF_X1 U280 ( .A(n246), .Z(n304) );
  NAND2_X1 U281 ( .A1(n320), .A2(n321), .ZN(n305) );
  AOI21_X1 U282 ( .B1(n338), .B2(n66), .A(n63), .ZN(n306) );
  AOI21_X1 U283 ( .B1(n338), .B2(n66), .A(n63), .ZN(n61) );
  BUF_X2 U284 ( .A(n227), .Z(n347) );
  XNOR2_X1 U285 ( .A(n245), .B(a[6]), .ZN(n307) );
  XNOR2_X1 U286 ( .A(n115), .B(n313), .ZN(n308) );
  NOR2_X1 U287 ( .A1(n125), .A2(n128), .ZN(n310) );
  OAI21_X1 U288 ( .B1(n301), .B2(n47), .A(n42), .ZN(n311) );
  OR2_X2 U289 ( .A1(n99), .A2(n102), .ZN(n337) );
  OAI21_X2 U290 ( .B1(n67), .B2(n69), .A(n68), .ZN(n66) );
  XNOR2_X1 U291 ( .A(n115), .B(n313), .ZN(n113) );
  XNOR2_X1 U292 ( .A(n120), .B(n117), .ZN(n313) );
  OAI21_X1 U293 ( .B1(n310), .B2(n306), .A(n60), .ZN(n314) );
  CLKBUF_X1 U294 ( .A(n71), .Z(n316) );
  CLKBUF_X1 U295 ( .A(n72), .Z(n317) );
  NAND2_X1 U296 ( .A1(n245), .A2(n319), .ZN(n320) );
  NAND2_X1 U297 ( .A1(n318), .A2(a[4]), .ZN(n321) );
  NAND2_X1 U298 ( .A1(n320), .A2(n321), .ZN(n229) );
  INV_X1 U299 ( .A(n245), .ZN(n318) );
  INV_X1 U300 ( .A(a[4]), .ZN(n319) );
  NAND2_X1 U301 ( .A1(n115), .A2(n120), .ZN(n322) );
  NAND2_X1 U302 ( .A1(n115), .A2(n117), .ZN(n323) );
  NAND2_X1 U303 ( .A1(n120), .A2(n117), .ZN(n324) );
  NAND3_X1 U304 ( .A1(n322), .A2(n323), .A3(n324), .ZN(n112) );
  NAND2_X1 U305 ( .A1(n305), .A2(n297), .ZN(n325) );
  NAND2_X1 U306 ( .A1(n229), .A2(n327), .ZN(n326) );
  OAI21_X1 U307 ( .B1(n331), .B2(n288), .A(n38), .ZN(n328) );
  OAI22_X1 U308 ( .A1(n234), .A2(n203), .B1(n202), .B2(n340), .ZN(n329) );
  INV_X1 U309 ( .A(n140), .ZN(n330) );
  BUF_X2 U310 ( .A(n238), .Z(n340) );
  AOI21_X1 U311 ( .B1(n50), .B2(n294), .A(n285), .ZN(n331) );
  AOI21_X1 U312 ( .B1(n50), .B2(n58), .A(n51), .ZN(n332) );
  AOI21_X1 U313 ( .B1(n315), .B2(n336), .A(n293), .ZN(n333) );
  XNOR2_X1 U314 ( .A(n48), .B(n5), .ZN(product[9]) );
  NAND2_X1 U315 ( .A1(n85), .A2(n47), .ZN(n5) );
  INV_X1 U316 ( .A(n46), .ZN(n85) );
  INV_X1 U317 ( .A(n47), .ZN(n45) );
  INV_X1 U318 ( .A(n311), .ZN(n38) );
  NAND2_X1 U319 ( .A1(n81), .A2(n21), .ZN(n1) );
  INV_X1 U320 ( .A(n20), .ZN(n81) );
  NAND2_X1 U321 ( .A1(n336), .A2(n30), .ZN(n2) );
  AOI21_X1 U322 ( .B1(n315), .B2(n336), .A(n293), .ZN(n26) );
  NOR2_X1 U323 ( .A1(n107), .A2(n112), .ZN(n46) );
  NAND2_X1 U324 ( .A1(n88), .A2(n60), .ZN(n8) );
  INV_X1 U325 ( .A(n310), .ZN(n88) );
  NAND2_X1 U326 ( .A1(n286), .A2(n42), .ZN(n4) );
  NAND2_X1 U327 ( .A1(n107), .A2(n112), .ZN(n47) );
  AOI21_X1 U328 ( .B1(n335), .B2(n78), .A(n75), .ZN(n73) );
  INV_X1 U329 ( .A(n77), .ZN(n75) );
  INV_X1 U330 ( .A(n80), .ZN(n78) );
  NAND2_X1 U331 ( .A1(n338), .A2(n65), .ZN(n9) );
  XOR2_X1 U332 ( .A(n57), .B(n7), .Z(product[7]) );
  NAND2_X1 U333 ( .A1(n87), .A2(n56), .ZN(n7) );
  INV_X1 U334 ( .A(n55), .ZN(n87) );
  XNOR2_X1 U335 ( .A(n12), .B(n78), .ZN(product[2]) );
  NAND2_X1 U336 ( .A1(n335), .A2(n77), .ZN(n12) );
  NAND2_X1 U337 ( .A1(n337), .A2(n35), .ZN(n3) );
  NOR2_X1 U338 ( .A1(n119), .A2(n124), .ZN(n55) );
  OR2_X1 U339 ( .A1(n169), .A2(n157), .ZN(n116) );
  NAND2_X1 U340 ( .A1(n91), .A2(n317), .ZN(n11) );
  INV_X1 U341 ( .A(n316), .ZN(n91) );
  INV_X1 U342 ( .A(n94), .ZN(n95) );
  NOR2_X1 U343 ( .A1(n96), .A2(n95), .ZN(n20) );
  OR2_X1 U344 ( .A1(n182), .A2(n175), .ZN(n335) );
  XOR2_X1 U345 ( .A(n10), .B(n69), .Z(product[4]) );
  NAND2_X1 U346 ( .A1(n90), .A2(n68), .ZN(n10) );
  INV_X1 U347 ( .A(n67), .ZN(n90) );
  NAND2_X1 U348 ( .A1(n119), .A2(n124), .ZN(n56) );
  NOR2_X1 U349 ( .A1(n125), .A2(n128), .ZN(n59) );
  XNOR2_X1 U350 ( .A(n54), .B(n6), .ZN(product[8]) );
  NAND2_X1 U351 ( .A1(n342), .A2(n53), .ZN(n6) );
  OAI21_X1 U352 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  OR2_X1 U353 ( .A1(n129), .A2(n132), .ZN(n338) );
  NAND2_X1 U354 ( .A1(n125), .A2(n128), .ZN(n60) );
  INV_X1 U355 ( .A(n70), .ZN(n69) );
  NAND2_X1 U356 ( .A1(n96), .A2(n95), .ZN(n21) );
  NAND2_X1 U357 ( .A1(n129), .A2(n132), .ZN(n65) );
  AND2_X1 U358 ( .A1(n347), .A2(n143), .ZN(n175) );
  INV_X1 U359 ( .A(n14), .ZN(product[15]) );
  AND2_X1 U360 ( .A1(n287), .A2(n80), .ZN(product[1]) );
  OR2_X1 U361 ( .A1(n347), .A2(n243), .ZN(n219) );
  AND2_X1 U362 ( .A1(n347), .A2(n140), .ZN(n167) );
  OR2_X1 U363 ( .A1(n347), .A2(n241), .ZN(n201) );
  NOR2_X1 U364 ( .A1(n133), .A2(n134), .ZN(n67) );
  INV_X1 U365 ( .A(n139), .ZN(n160) );
  INV_X1 U366 ( .A(n100), .ZN(n101) );
  AND2_X1 U367 ( .A1(n347), .A2(n137), .ZN(n159) );
  INV_X1 U368 ( .A(n136), .ZN(n152) );
  NAND2_X1 U369 ( .A1(n133), .A2(n134), .ZN(n68) );
  OR2_X1 U370 ( .A1(n347), .A2(n240), .ZN(n192) );
  OR2_X1 U371 ( .A1(n347), .A2(n242), .ZN(n210) );
  INV_X1 U372 ( .A(n146), .ZN(n255) );
  NAND2_X1 U373 ( .A1(n228), .A2(n307), .ZN(n232) );
  AND2_X1 U374 ( .A1(n347), .A2(n146), .ZN(product[0]) );
  NAND2_X1 U375 ( .A1(n135), .A2(n150), .ZN(n72) );
  OAI21_X1 U376 ( .B1(n301), .B2(n47), .A(n42), .ZN(n40) );
  NOR2_X1 U377 ( .A1(n46), .A2(n41), .ZN(n39) );
  OAI22_X1 U378 ( .A1(n292), .A2(n214), .B1(n213), .B2(n255), .ZN(n179) );
  OAI22_X1 U379 ( .A1(n292), .A2(n215), .B1(n214), .B2(n255), .ZN(n180) );
  OAI22_X1 U380 ( .A1(n235), .A2(n213), .B1(n212), .B2(n255), .ZN(n178) );
  OAI22_X1 U381 ( .A1(n235), .A2(n212), .B1(n211), .B2(n255), .ZN(n177) );
  OAI22_X1 U382 ( .A1(n290), .A2(n292), .B1(n290), .B2(n255), .ZN(n145) );
  OAI22_X1 U383 ( .A1(n292), .A2(n216), .B1(n215), .B2(n255), .ZN(n181) );
  OAI22_X1 U384 ( .A1(n292), .A2(n243), .B1(n219), .B2(n255), .ZN(n151) );
  OAI22_X1 U385 ( .A1(n292), .A2(n218), .B1(n217), .B2(n255), .ZN(n183) );
  XNOR2_X1 U386 ( .A(n245), .B(a[6]), .ZN(n236) );
  XNOR2_X1 U387 ( .A(n247), .B(a[2]), .ZN(n238) );
  XNOR2_X1 U388 ( .A(n347), .B(n244), .ZN(n191) );
  XNOR2_X1 U389 ( .A(n244), .B(b[4]), .ZN(n187) );
  XNOR2_X1 U390 ( .A(n244), .B(b[5]), .ZN(n186) );
  XNOR2_X1 U391 ( .A(n244), .B(b[6]), .ZN(n185) );
  INV_X1 U392 ( .A(n244), .ZN(n240) );
  XOR2_X1 U393 ( .A(n244), .B(a[6]), .Z(n228) );
  NAND2_X1 U394 ( .A1(n230), .A2(n238), .ZN(n341) );
  NAND2_X1 U395 ( .A1(n230), .A2(n238), .ZN(n234) );
  OR2_X1 U396 ( .A1(n308), .A2(n118), .ZN(n342) );
  NAND2_X1 U397 ( .A1(n229), .A2(n237), .ZN(n344) );
  NAND2_X1 U398 ( .A1(n305), .A2(n298), .ZN(n345) );
  NAND2_X1 U399 ( .A1(n305), .A2(n237), .ZN(n233) );
  XNOR2_X1 U400 ( .A(n246), .B(a[4]), .ZN(n237) );
  XOR2_X1 U401 ( .A(n8), .B(n306), .Z(product[6]) );
  INV_X1 U402 ( .A(n145), .ZN(n176) );
  INV_X1 U403 ( .A(n110), .ZN(n111) );
  NAND2_X1 U404 ( .A1(n103), .A2(n106), .ZN(n42) );
  XNOR2_X1 U405 ( .A(n9), .B(n66), .ZN(product[5]) );
  NAND2_X1 U406 ( .A1(n182), .A2(n175), .ZN(n77) );
  OAI22_X1 U407 ( .A1(n292), .A2(n217), .B1(n216), .B2(n255), .ZN(n182) );
  INV_X1 U408 ( .A(n142), .ZN(n168) );
  INV_X1 U409 ( .A(n314), .ZN(n57) );
  NOR2_X1 U410 ( .A1(n135), .A2(n150), .ZN(n71) );
  OAI22_X1 U411 ( .A1(n184), .A2(n334), .B1(n184), .B2(n343), .ZN(n136) );
  OAI22_X1 U412 ( .A1(n334), .A2(n185), .B1(n184), .B2(n343), .ZN(n94) );
  OAI22_X1 U413 ( .A1(n334), .A2(n188), .B1(n187), .B2(n343), .ZN(n155) );
  OAI22_X1 U414 ( .A1(n334), .A2(n187), .B1(n186), .B2(n343), .ZN(n154) );
  OAI22_X1 U415 ( .A1(n334), .A2(n186), .B1(n185), .B2(n343), .ZN(n153) );
  OAI22_X1 U416 ( .A1(n334), .A2(n190), .B1(n189), .B2(n236), .ZN(n157) );
  INV_X1 U417 ( .A(n236), .ZN(n137) );
  OAI22_X1 U418 ( .A1(n334), .A2(n189), .B1(n188), .B2(n236), .ZN(n156) );
  OAI22_X1 U419 ( .A1(n232), .A2(n240), .B1(n192), .B2(n236), .ZN(n148) );
  OAI22_X1 U420 ( .A1(n232), .A2(n191), .B1(n190), .B2(n236), .ZN(n158) );
  XNOR2_X1 U421 ( .A(n300), .B(b[4]), .ZN(n196) );
  XNOR2_X1 U422 ( .A(n291), .B(b[5]), .ZN(n195) );
  XNOR2_X1 U423 ( .A(n291), .B(b[6]), .ZN(n194) );
  XNOR2_X1 U424 ( .A(n347), .B(n300), .ZN(n200) );
  INV_X1 U425 ( .A(n245), .ZN(n241) );
  NOR2_X1 U426 ( .A1(n52), .A2(n55), .ZN(n50) );
  NOR2_X1 U427 ( .A1(n113), .A2(n118), .ZN(n52) );
  NAND2_X1 U428 ( .A1(n308), .A2(n118), .ZN(n53) );
  CLKBUF_X1 U429 ( .A(n328), .Z(n346) );
  OAI21_X1 U430 ( .B1(n331), .B2(n288), .A(n38), .ZN(n36) );
  INV_X1 U431 ( .A(n333), .ZN(n24) );
  OAI21_X1 U432 ( .B1(n26), .B2(n20), .A(n21), .ZN(n19) );
  XNOR2_X1 U433 ( .A(n309), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U434 ( .A(n309), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U435 ( .A(n309), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U436 ( .A(n347), .B(n309), .ZN(n218) );
  INV_X1 U437 ( .A(n65), .ZN(n63) );
  AOI21_X1 U438 ( .B1(n50), .B2(n314), .A(n285), .ZN(n49) );
  OAI21_X1 U439 ( .B1(n59), .B2(n61), .A(n60), .ZN(n58) );
  XOR2_X1 U440 ( .A(n43), .B(n4), .Z(product[10]) );
  XOR2_X1 U441 ( .A(n31), .B(n2), .Z(product[12]) );
  XOR2_X1 U442 ( .A(n11), .B(n73), .Z(product[3]) );
  OAI21_X1 U443 ( .B1(n71), .B2(n73), .A(n72), .ZN(n70) );
  NAND2_X1 U444 ( .A1(n183), .A2(n151), .ZN(n80) );
  NOR2_X1 U445 ( .A1(n25), .A2(n20), .ZN(n18) );
  NAND2_X1 U446 ( .A1(n337), .A2(n336), .ZN(n25) );
  NAND2_X1 U447 ( .A1(n39), .A2(n302), .ZN(n16) );
  AOI21_X1 U448 ( .B1(n40), .B2(n18), .A(n19), .ZN(n17) );
  OAI21_X1 U449 ( .B1(n52), .B2(n56), .A(n53), .ZN(n51) );
  XOR2_X1 U450 ( .A(n22), .B(n1), .Z(product[13]) );
  OAI22_X1 U451 ( .A1(n344), .A2(n199), .B1(n198), .B2(n330), .ZN(n165) );
  OAI22_X1 U452 ( .A1(n326), .A2(n198), .B1(n197), .B2(n298), .ZN(n164) );
  OAI22_X1 U453 ( .A1(n345), .A2(n197), .B1(n196), .B2(n297), .ZN(n163) );
  OAI22_X1 U454 ( .A1(n344), .A2(n194), .B1(n193), .B2(n330), .ZN(n100) );
  OAI22_X1 U455 ( .A1(n344), .A2(n196), .B1(n195), .B2(n297), .ZN(n162) );
  INV_X1 U456 ( .A(n298), .ZN(n140) );
  OAI22_X1 U457 ( .A1(n193), .A2(n344), .B1(n193), .B2(n330), .ZN(n139) );
  OAI22_X1 U458 ( .A1(n325), .A2(n195), .B1(n194), .B2(n298), .ZN(n161) );
  XNOR2_X1 U459 ( .A(n312), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U460 ( .A(n312), .B(b[5]), .ZN(n204) );
  OAI22_X1 U461 ( .A1(n233), .A2(n241), .B1(n201), .B2(n297), .ZN(n149) );
  OAI22_X1 U462 ( .A1(n233), .A2(n200), .B1(n199), .B2(n298), .ZN(n166) );
  INV_X1 U463 ( .A(n312), .ZN(n242) );
  XNOR2_X1 U464 ( .A(n312), .B(b[6]), .ZN(n203) );
  XNOR2_X1 U465 ( .A(n347), .B(n312), .ZN(n209) );
  XOR2_X1 U466 ( .A(n246), .B(a[2]), .Z(n230) );
  XOR2_X1 U467 ( .A(n247), .B(n146), .Z(n231) );
  INV_X1 U468 ( .A(n309), .ZN(n243) );
  XNOR2_X1 U469 ( .A(n244), .B(b[7]), .ZN(n184) );
  XNOR2_X1 U470 ( .A(n300), .B(b[7]), .ZN(n193) );
  XNOR2_X1 U471 ( .A(n309), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U472 ( .A(n304), .B(b[7]), .ZN(n202) );
  XNOR2_X1 U473 ( .A(n312), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U474 ( .A(n289), .B(b[3]), .ZN(n197) );
  XNOR2_X1 U475 ( .A(n244), .B(b[3]), .ZN(n188) );
  XNOR2_X1 U476 ( .A(n309), .B(b[3]), .ZN(n215) );
  AOI21_X1 U477 ( .B1(n48), .B2(n85), .A(n45), .ZN(n43) );
  XNOR2_X1 U478 ( .A(n244), .B(b[2]), .ZN(n189) );
  XNOR2_X1 U479 ( .A(n312), .B(b[2]), .ZN(n207) );
  XNOR2_X1 U480 ( .A(n289), .B(b[2]), .ZN(n198) );
  XNOR2_X1 U481 ( .A(n309), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U482 ( .A(n244), .B(b[1]), .ZN(n190) );
  XNOR2_X1 U483 ( .A(n291), .B(b[1]), .ZN(n199) );
  XNOR2_X1 U484 ( .A(n312), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U485 ( .A(n309), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U486 ( .A(n346), .B(n3), .ZN(product[11]) );
  AOI21_X1 U487 ( .B1(n328), .B2(n337), .A(n295), .ZN(n31) );
  AOI21_X1 U488 ( .B1(n36), .B2(n296), .A(n24), .ZN(n22) );
  OAI21_X1 U489 ( .B1(n332), .B2(n16), .A(n17), .ZN(n15) );
  INV_X1 U490 ( .A(n49), .ZN(n48) );
  OAI22_X1 U491 ( .A1(n234), .A2(n204), .B1(n203), .B2(n340), .ZN(n169) );
  OAI22_X1 U492 ( .A1(n234), .A2(n207), .B1(n206), .B2(n340), .ZN(n172) );
  OAI22_X1 U493 ( .A1(n234), .A2(n206), .B1(n205), .B2(n340), .ZN(n171) );
  OAI22_X1 U494 ( .A1(n205), .A2(n341), .B1(n204), .B2(n340), .ZN(n170) );
  OAI22_X1 U495 ( .A1(n234), .A2(n208), .B1(n207), .B2(n340), .ZN(n173) );
  OAI22_X1 U496 ( .A1(n234), .A2(n242), .B1(n210), .B2(n340), .ZN(n150) );
  OAI22_X1 U497 ( .A1(n341), .A2(n203), .B1(n202), .B2(n340), .ZN(n110) );
  OAI22_X1 U498 ( .A1(n341), .A2(n202), .B1(n202), .B2(n340), .ZN(n142) );
  INV_X1 U499 ( .A(n340), .ZN(n143) );
  OAI22_X1 U500 ( .A1(n299), .A2(n209), .B1(n208), .B2(n340), .ZN(n174) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1 ( clk, ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;
  input clk;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1_DW_mult_tc_1 mult_57 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module add_layer_WIDTH16_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  AND2_X1 U106 ( .A1(n157), .A2(n71), .ZN(SUM[0]) );
  CLKBUF_X1 U107 ( .A(n38), .Z(n143) );
  CLKBUF_X1 U108 ( .A(n35), .Z(n144) );
  CLKBUF_X1 U109 ( .A(n67), .Z(n145) );
  AOI21_X1 U110 ( .B1(n144), .B2(n153), .A(n32), .ZN(n146) );
  AOI21_X1 U111 ( .B1(n145), .B2(n150), .A(n64), .ZN(n147) );
  CLKBUF_X1 U112 ( .A(n54), .Z(n148) );
  XNOR2_X1 U113 ( .A(n16), .B(n149), .ZN(SUM[15]) );
  XOR2_X1 U114 ( .A(B[15]), .B(A[15]), .Z(n149) );
  INV_X1 U115 ( .A(n34), .ZN(n32) );
  INV_X1 U116 ( .A(n58), .ZN(n56) );
  INV_X1 U117 ( .A(n50), .ZN(n48) );
  OAI21_X1 U118 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  AOI21_X1 U119 ( .B1(n43), .B2(n155), .A(n40), .ZN(n38) );
  INV_X1 U120 ( .A(n42), .ZN(n40) );
  AOI21_X1 U121 ( .B1(n67), .B2(n150), .A(n64), .ZN(n62) );
  INV_X1 U122 ( .A(n66), .ZN(n64) );
  NAND2_X1 U123 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U124 ( .A(n28), .ZN(n76) );
  NAND2_X1 U125 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U126 ( .A(n52), .ZN(n82) );
  NAND2_X1 U127 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U128 ( .A(n44), .ZN(n80) );
  NAND2_X1 U129 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U130 ( .A(n36), .ZN(n78) );
  NAND2_X1 U131 ( .A1(n155), .A2(n42), .ZN(n7) );
  NAND2_X1 U132 ( .A1(n156), .A2(n20), .ZN(n2) );
  NAND2_X1 U133 ( .A1(n154), .A2(n26), .ZN(n3) );
  NAND2_X1 U134 ( .A1(n151), .A2(n50), .ZN(n9) );
  NAND2_X1 U135 ( .A1(n153), .A2(n34), .ZN(n5) );
  NAND2_X1 U136 ( .A1(n152), .A2(n58), .ZN(n11) );
  XNOR2_X1 U137 ( .A(n145), .B(n13), .ZN(SUM[2]) );
  NAND2_X1 U138 ( .A1(n150), .A2(n66), .ZN(n13) );
  NAND2_X1 U139 ( .A1(n86), .A2(n69), .ZN(n14) );
  INV_X1 U140 ( .A(n68), .ZN(n86) );
  NAND2_X1 U141 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U142 ( .A(n60), .ZN(n84) );
  INV_X1 U143 ( .A(n20), .ZN(n18) );
  NOR2_X1 U144 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  INV_X1 U145 ( .A(n26), .ZN(n24) );
  OR2_X1 U146 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  NOR2_X1 U147 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  NOR2_X1 U148 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NOR2_X1 U151 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NAND2_X1 U152 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U153 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U154 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U155 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U156 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  OR2_X1 U157 ( .A1(A[6]), .A2(B[6]), .ZN(n151) );
  OR2_X1 U158 ( .A1(A[4]), .A2(B[4]), .ZN(n152) );
  OR2_X1 U159 ( .A1(A[10]), .A2(B[10]), .ZN(n153) );
  OR2_X1 U160 ( .A1(A[12]), .A2(B[12]), .ZN(n154) );
  OR2_X1 U161 ( .A1(A[8]), .A2(B[8]), .ZN(n155) );
  NAND2_X1 U162 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U163 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U164 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  NAND2_X1 U165 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U166 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  OR2_X1 U167 ( .A1(A[14]), .A2(B[14]), .ZN(n156) );
  NAND2_X1 U168 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  OR2_X1 U169 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  NAND2_X1 U170 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  XOR2_X1 U171 ( .A(n14), .B(n71), .Z(SUM[1]) );
  AOI21_X1 U172 ( .B1(n51), .B2(n151), .A(n48), .ZN(n46) );
  NAND2_X1 U173 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  OAI21_X1 U174 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  AOI21_X1 U175 ( .B1(n59), .B2(n152), .A(n56), .ZN(n54) );
  OAI21_X1 U176 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  XOR2_X1 U177 ( .A(n147), .B(n12), .Z(SUM[3]) );
  XNOR2_X1 U178 ( .A(n43), .B(n7), .ZN(SUM[8]) );
  OAI21_X1 U179 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  XOR2_X1 U180 ( .A(n146), .B(n4), .Z(SUM[11]) );
  AOI21_X1 U181 ( .B1(n35), .B2(n153), .A(n32), .ZN(n30) );
  OAI21_X1 U182 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  XOR2_X1 U183 ( .A(n46), .B(n8), .Z(SUM[7]) );
  XNOR2_X1 U184 ( .A(n27), .B(n3), .ZN(SUM[12]) );
  XNOR2_X1 U185 ( .A(n144), .B(n5), .ZN(SUM[10]) );
  XNOR2_X1 U186 ( .A(n51), .B(n9), .ZN(SUM[6]) );
  XOR2_X1 U187 ( .A(n143), .B(n6), .Z(SUM[9]) );
  OAI21_X1 U188 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  XOR2_X1 U189 ( .A(n148), .B(n10), .Z(SUM[5]) );
  XNOR2_X1 U190 ( .A(n59), .B(n11), .ZN(SUM[4]) );
  XNOR2_X1 U191 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  AOI21_X1 U192 ( .B1(n21), .B2(n156), .A(n18), .ZN(n16) );
  INV_X1 U193 ( .A(n22), .ZN(n73) );
  NAND2_X1 U194 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  AOI21_X1 U195 ( .B1(n154), .B2(n27), .A(n24), .ZN(n22) );
endmodule


module add_layer_WIDTH16_6 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_6_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n36, n37,
         n38, n40, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n56,
         n58, n59, n60, n61, n62, n64, n66, n67, n68, n69, n71, n73, n76, n78,
         n80, n82, n84, n86, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156;

  FA_X1 U12 ( .A(A[13]), .B(B[13]), .CI(n73), .CO(n21), .S(SUM[13]) );
  OR2_X1 U106 ( .A1(A[0]), .A2(B[0]), .ZN(n142) );
  CLKBUF_X1 U107 ( .A(n38), .Z(n143) );
  CLKBUF_X1 U108 ( .A(n35), .Z(n144) );
  CLKBUF_X1 U109 ( .A(n67), .Z(n145) );
  AOI21_X1 U110 ( .B1(n144), .B2(n153), .A(n32), .ZN(n146) );
  AOI21_X1 U111 ( .B1(n145), .B2(n156), .A(n64), .ZN(n147) );
  CLKBUF_X1 U112 ( .A(n54), .Z(n148) );
  XNOR2_X1 U113 ( .A(n16), .B(n149), .ZN(SUM[15]) );
  XOR2_X1 U114 ( .A(B[15]), .B(A[15]), .Z(n149) );
  INV_X1 U115 ( .A(n42), .ZN(n40) );
  INV_X1 U116 ( .A(n34), .ZN(n32) );
  INV_X1 U117 ( .A(n50), .ZN(n48) );
  AOI21_X1 U118 ( .B1(n67), .B2(n156), .A(n64), .ZN(n62) );
  INV_X1 U119 ( .A(n66), .ZN(n64) );
  OAI21_X1 U120 ( .B1(n62), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X1 U121 ( .B1(n59), .B2(n150), .A(n56), .ZN(n54) );
  INV_X1 U122 ( .A(n58), .ZN(n56) );
  NAND2_X1 U123 ( .A1(n76), .A2(n29), .ZN(n4) );
  INV_X1 U124 ( .A(n28), .ZN(n76) );
  NAND2_X1 U125 ( .A1(n84), .A2(n61), .ZN(n12) );
  INV_X1 U126 ( .A(n60), .ZN(n84) );
  NAND2_X1 U127 ( .A1(n82), .A2(n53), .ZN(n10) );
  INV_X1 U128 ( .A(n52), .ZN(n82) );
  NAND2_X1 U129 ( .A1(n80), .A2(n45), .ZN(n8) );
  INV_X1 U130 ( .A(n44), .ZN(n80) );
  NAND2_X1 U131 ( .A1(n78), .A2(n37), .ZN(n6) );
  INV_X1 U132 ( .A(n36), .ZN(n78) );
  NAND2_X1 U133 ( .A1(n153), .A2(n34), .ZN(n5) );
  NAND2_X1 U134 ( .A1(n154), .A2(n26), .ZN(n3) );
  NAND2_X1 U135 ( .A1(n151), .A2(n42), .ZN(n7) );
  NAND2_X1 U136 ( .A1(n150), .A2(n58), .ZN(n11) );
  NAND2_X1 U137 ( .A1(n152), .A2(n50), .ZN(n9) );
  XOR2_X1 U138 ( .A(n14), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U139 ( .A1(n86), .A2(n69), .ZN(n14) );
  XNOR2_X1 U140 ( .A(n21), .B(n2), .ZN(SUM[14]) );
  NAND2_X1 U141 ( .A1(n155), .A2(n20), .ZN(n2) );
  INV_X1 U142 ( .A(n20), .ZN(n18) );
  NAND2_X1 U143 ( .A1(A[0]), .A2(B[0]), .ZN(n71) );
  INV_X1 U144 ( .A(n26), .ZN(n24) );
  NOR2_X1 U145 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  NOR2_X1 U146 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  OR2_X1 U147 ( .A1(A[4]), .A2(B[4]), .ZN(n150) );
  NOR2_X1 U148 ( .A1(A[5]), .A2(B[5]), .ZN(n52) );
  NOR2_X1 U149 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(B[9]), .ZN(n36) );
  NOR2_X1 U151 ( .A1(A[11]), .A2(B[11]), .ZN(n28) );
  NAND2_X1 U152 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U153 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U154 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U155 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U156 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U157 ( .A1(A[14]), .A2(B[14]), .ZN(n20) );
  NAND2_X1 U158 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  OR2_X1 U159 ( .A1(A[8]), .A2(B[8]), .ZN(n151) );
  OR2_X1 U160 ( .A1(A[6]), .A2(B[6]), .ZN(n152) );
  OR2_X1 U161 ( .A1(A[10]), .A2(B[10]), .ZN(n153) );
  OR2_X1 U162 ( .A1(A[12]), .A2(B[12]), .ZN(n154) );
  OR2_X1 U163 ( .A1(A[14]), .A2(B[14]), .ZN(n155) );
  NAND2_X1 U164 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U165 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U166 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U167 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  OR2_X1 U168 ( .A1(A[2]), .A2(B[2]), .ZN(n156) );
  AND2_X1 U169 ( .A1(n142), .A2(n71), .ZN(SUM[0]) );
  XNOR2_X1 U170 ( .A(n145), .B(n13), .ZN(SUM[2]) );
  OAI21_X1 U171 ( .B1(n68), .B2(n71), .A(n69), .ZN(n67) );
  AOI21_X1 U172 ( .B1(n51), .B2(n152), .A(n48), .ZN(n46) );
  OAI21_X1 U173 ( .B1(n46), .B2(n44), .A(n45), .ZN(n43) );
  NAND2_X1 U174 ( .A1(n156), .A2(n66), .ZN(n13) );
  NAND2_X1 U175 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  XNOR2_X1 U176 ( .A(n43), .B(n7), .ZN(SUM[8]) );
  INV_X1 U177 ( .A(n68), .ZN(n86) );
  AOI21_X1 U178 ( .B1(n43), .B2(n151), .A(n40), .ZN(n38) );
  OAI21_X1 U179 ( .B1(n54), .B2(n52), .A(n53), .ZN(n51) );
  XNOR2_X1 U180 ( .A(n51), .B(n9), .ZN(SUM[6]) );
  XOR2_X1 U181 ( .A(n46), .B(n8), .Z(SUM[7]) );
  XNOR2_X1 U182 ( .A(n144), .B(n5), .ZN(SUM[10]) );
  XOR2_X1 U183 ( .A(n148), .B(n10), .Z(SUM[5]) );
  AOI21_X1 U184 ( .B1(n35), .B2(n153), .A(n32), .ZN(n30) );
  OAI21_X1 U185 ( .B1(n38), .B2(n36), .A(n37), .ZN(n35) );
  XNOR2_X1 U186 ( .A(n59), .B(n11), .ZN(SUM[4]) );
  XOR2_X1 U187 ( .A(n143), .B(n6), .Z(SUM[9]) );
  INV_X1 U188 ( .A(n22), .ZN(n73) );
  XNOR2_X1 U189 ( .A(n27), .B(n3), .ZN(SUM[12]) );
  XOR2_X1 U190 ( .A(n147), .B(n12), .Z(SUM[3]) );
  AOI21_X1 U191 ( .B1(n154), .B2(n27), .A(n24), .ZN(n22) );
  OAI21_X1 U192 ( .B1(n30), .B2(n28), .A(n29), .ZN(n27) );
  NAND2_X1 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  AOI21_X1 U194 ( .B1(n21), .B2(n155), .A(n18), .ZN(n16) );
  XOR2_X1 U195 ( .A(n146), .B(n4), .Z(SUM[11]) );
endmodule


module add_layer_WIDTH16_5 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_5_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module add_layer_WIDTH16_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37,
         n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70,
         n71, n73, n75, n77, n79, n81, n82, n83, n84, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n71), .CO(n16), .S(SUM[14]) );
  NAND2_X1 U104 ( .A1(A[2]), .A2(B[2]), .ZN(n64) );
  AND2_X1 U105 ( .A1(n157), .A2(n70), .ZN(SUM[0]) );
  CLKBUF_X1 U106 ( .A(n46), .Z(n141) );
  AOI21_X1 U107 ( .B1(n141), .B2(n156), .A(n43), .ZN(n142) );
  CLKBUF_X1 U108 ( .A(n30), .Z(n143) );
  AOI21_X1 U109 ( .B1(n143), .B2(n154), .A(n27), .ZN(n144) );
  CLKBUF_X1 U110 ( .A(n54), .Z(n145) );
  CLKBUF_X1 U111 ( .A(n38), .Z(n146) );
  CLKBUF_X1 U112 ( .A(n57), .Z(n147) );
  AOI21_X1 U113 ( .B1(n54), .B2(n152), .A(n51), .ZN(n148) );
  AOI21_X1 U114 ( .B1(n38), .B2(n153), .A(n35), .ZN(n149) );
  NOR2_X1 U115 ( .A1(A[3]), .A2(B[3]), .ZN(n150) );
  OR2_X1 U116 ( .A1(A[5]), .A2(B[5]), .ZN(n152) );
  INV_X1 U117 ( .A(n37), .ZN(n35) );
  INV_X1 U118 ( .A(n29), .ZN(n27) );
  AOI21_X1 U119 ( .B1(n145), .B2(n152), .A(n51), .ZN(n49) );
  INV_X1 U120 ( .A(n53), .ZN(n51) );
  OAI21_X1 U121 ( .B1(n148), .B2(n47), .A(n48), .ZN(n46) );
  AOI21_X1 U122 ( .B1(n66), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U123 ( .B1(n46), .B2(n156), .A(n43), .ZN(n41) );
  INV_X1 U124 ( .A(n45), .ZN(n43) );
  NAND2_X1 U125 ( .A1(n73), .A2(n24), .ZN(n3) );
  INV_X1 U126 ( .A(n23), .ZN(n73) );
  NAND2_X1 U127 ( .A1(n154), .A2(n29), .ZN(n4) );
  NAND2_X1 U128 ( .A1(n155), .A2(n21), .ZN(n2) );
  NAND2_X1 U129 ( .A1(n84), .A2(n68), .ZN(n14) );
  INV_X1 U130 ( .A(n67), .ZN(n84) );
  OAI21_X1 U131 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  XNOR2_X1 U132 ( .A(n145), .B(n10), .ZN(SUM[5]) );
  NAND2_X1 U133 ( .A1(n152), .A2(n53), .ZN(n10) );
  NAND2_X1 U134 ( .A1(n83), .A2(n64), .ZN(n13) );
  INV_X1 U135 ( .A(n63), .ZN(n83) );
  NAND2_X1 U136 ( .A1(n82), .A2(n61), .ZN(n12) );
  NAND2_X1 U137 ( .A1(n156), .A2(n45), .ZN(n8) );
  NAND2_X1 U138 ( .A1(n153), .A2(n37), .ZN(n6) );
  NAND2_X1 U139 ( .A1(n79), .A2(n48), .ZN(n9) );
  INV_X1 U140 ( .A(n47), .ZN(n79) );
  NAND2_X1 U141 ( .A1(n77), .A2(n40), .ZN(n7) );
  INV_X1 U142 ( .A(n39), .ZN(n77) );
  NAND2_X1 U143 ( .A1(n75), .A2(n32), .ZN(n5) );
  INV_X1 U144 ( .A(n31), .ZN(n75) );
  NAND2_X1 U145 ( .A1(n81), .A2(n56), .ZN(n11) );
  INV_X1 U146 ( .A(n55), .ZN(n81) );
  XNOR2_X1 U147 ( .A(n16), .B(n151), .ZN(SUM[15]) );
  XNOR2_X1 U148 ( .A(B[15]), .B(A[15]), .ZN(n151) );
  NOR2_X1 U149 ( .A1(A[6]), .A2(B[6]), .ZN(n47) );
  NOR2_X1 U150 ( .A1(A[8]), .A2(B[8]), .ZN(n39) );
  NOR2_X1 U151 ( .A1(A[4]), .A2(B[4]), .ZN(n55) );
  NOR2_X1 U152 ( .A1(A[10]), .A2(B[10]), .ZN(n31) );
  NOR2_X1 U153 ( .A1(A[12]), .A2(B[12]), .ZN(n23) );
  INV_X1 U154 ( .A(n21), .ZN(n19) );
  NAND2_X1 U155 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U156 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U157 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U158 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U159 ( .A1(A[13]), .A2(B[13]), .ZN(n21) );
  NAND2_X1 U160 ( .A1(A[6]), .A2(B[6]), .ZN(n48) );
  OR2_X1 U161 ( .A1(A[9]), .A2(B[9]), .ZN(n153) );
  OR2_X1 U162 ( .A1(A[11]), .A2(B[11]), .ZN(n154) );
  OR2_X1 U163 ( .A1(A[13]), .A2(B[13]), .ZN(n155) );
  OR2_X1 U164 ( .A1(A[7]), .A2(B[7]), .ZN(n156) );
  NAND2_X1 U165 ( .A1(A[8]), .A2(B[8]), .ZN(n40) );
  NAND2_X1 U166 ( .A1(A[4]), .A2(B[4]), .ZN(n56) );
  NAND2_X1 U167 ( .A1(A[10]), .A2(B[10]), .ZN(n32) );
  NAND2_X1 U168 ( .A1(A[12]), .A2(B[12]), .ZN(n24) );
  XNOR2_X1 U169 ( .A(n62), .B(n12), .ZN(SUM[3]) );
  XOR2_X1 U170 ( .A(n65), .B(n13), .Z(SUM[2]) );
  OR2_X1 U171 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  NOR2_X2 U172 ( .A1(A[2]), .A2(B[2]), .ZN(n63) );
  XNOR2_X1 U173 ( .A(n146), .B(n6), .ZN(SUM[9]) );
  XOR2_X1 U174 ( .A(n14), .B(n70), .Z(SUM[1]) );
  AOI21_X1 U175 ( .B1(n146), .B2(n153), .A(n35), .ZN(n33) );
  OAI21_X1 U176 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  NAND2_X1 U177 ( .A1(A[0]), .A2(B[0]), .ZN(n70) );
  NOR2_X1 U178 ( .A1(A[1]), .A2(B[1]), .ZN(n67) );
  NAND2_X1 U179 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  XOR2_X1 U180 ( .A(n142), .B(n7), .Z(SUM[8]) );
  XNOR2_X1 U181 ( .A(n143), .B(n4), .ZN(SUM[11]) );
  XNOR2_X1 U182 ( .A(n141), .B(n8), .ZN(SUM[7]) );
  XOR2_X1 U183 ( .A(n33), .B(n5), .Z(SUM[10]) );
  OAI21_X1 U184 ( .B1(n149), .B2(n31), .A(n32), .ZN(n30) );
  XOR2_X1 U185 ( .A(n49), .B(n9), .Z(SUM[6]) );
  OAI21_X1 U186 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  INV_X1 U187 ( .A(n66), .ZN(n65) );
  INV_X1 U188 ( .A(n17), .ZN(n71) );
  AOI21_X1 U189 ( .B1(n155), .B2(n22), .A(n19), .ZN(n17) );
  XNOR2_X1 U190 ( .A(n22), .B(n2), .ZN(SUM[13]) );
  XOR2_X1 U191 ( .A(n144), .B(n3), .Z(SUM[12]) );
  OAI21_X1 U192 ( .B1(n25), .B2(n23), .A(n24), .ZN(n22) );
  AOI21_X1 U193 ( .B1(n30), .B2(n154), .A(n27), .ZN(n25) );
  XOR2_X1 U194 ( .A(n147), .B(n11), .Z(SUM[4]) );
  OAI21_X1 U195 ( .B1(n67), .B2(n70), .A(n68), .ZN(n66) );
  NOR2_X1 U196 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NAND2_X1 U197 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
  OAI21_X1 U198 ( .B1(n60), .B2(n64), .A(n61), .ZN(n59) );
  NOR2_X1 U199 ( .A1(n63), .A2(n150), .ZN(n58) );
  INV_X1 U200 ( .A(n150), .ZN(n82) );
endmodule


module add_layer_WIDTH16_1 ( clk, a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [15:0] out;
  input clk;


  add_layer_WIDTH16_1_DW01_add_1 add_68 ( .A(a), .B(b), .CI(1'b0), .SUM(out)
         );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_1 ( clk, .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input clk, \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;
  wire   \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ;

  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_1 \genblk2.add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_1 ( clk, .in({
        \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , 
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , 
        \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , 
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] 
        }), out );
  output [15:0] out;
  input clk, \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] ,
         \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] ,
         \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] ,
         \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] ,
         \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] ,
         \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] ,
         \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] ,
         \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] ,
         \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] ,
         \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] ,
         \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] ,
         \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] ,
         \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] ,
         \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] ,
         \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] ,
         \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] ,
         \genblk2.inter[1][15] , \genblk2.inter[1][14] ,
         \genblk2.inter[1][13] , \genblk2.inter[1][12] ,
         \genblk2.inter[1][11] , \genblk2.inter[1][10] , \genblk2.inter[1][9] ,
         \genblk2.inter[1][8] , \genblk2.inter[1][7] , \genblk2.inter[1][6] ,
         \genblk2.inter[1][5] , \genblk2.inter[1][4] , \genblk2.inter[1][3] ,
         \genblk2.inter[1][2] , \genblk2.inter[1][1] , \genblk2.inter[1][0] ,
         \genblk2.inter[0][15] , \genblk2.inter[0][14] ,
         \genblk2.inter[0][13] , \genblk2.inter[0][12] ,
         \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] ,
         \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] ,
         \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] ,
         \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] ;

  DFF_X1 \add_in_reg[3][15]  ( .D(\in[3][15] ), .CK(clk), .Q(\add_in[3][15] )
         );
  DFF_X1 \add_in_reg[3][14]  ( .D(\in[3][14] ), .CK(clk), .Q(\add_in[3][14] )
         );
  DFF_X1 \add_in_reg[3][13]  ( .D(\in[3][13] ), .CK(clk), .Q(\add_in[3][13] )
         );
  DFF_X1 \add_in_reg[3][12]  ( .D(\in[3][12] ), .CK(clk), .Q(\add_in[3][12] )
         );
  DFF_X1 \add_in_reg[3][11]  ( .D(\in[3][11] ), .CK(clk), .Q(\add_in[3][11] )
         );
  DFF_X1 \add_in_reg[3][10]  ( .D(\in[3][10] ), .CK(clk), .Q(\add_in[3][10] )
         );
  DFF_X1 \add_in_reg[3][9]  ( .D(\in[3][9] ), .CK(clk), .Q(\add_in[3][9] ) );
  DFF_X1 \add_in_reg[3][8]  ( .D(\in[3][8] ), .CK(clk), .Q(\add_in[3][8] ) );
  DFF_X1 \add_in_reg[3][7]  ( .D(\in[3][7] ), .CK(clk), .Q(\add_in[3][7] ) );
  DFF_X1 \add_in_reg[3][6]  ( .D(\in[3][6] ), .CK(clk), .Q(\add_in[3][6] ) );
  DFF_X1 \add_in_reg[3][5]  ( .D(\in[3][5] ), .CK(clk), .Q(\add_in[3][5] ) );
  DFF_X1 \add_in_reg[3][4]  ( .D(\in[3][4] ), .CK(clk), .Q(\add_in[3][4] ) );
  DFF_X1 \add_in_reg[3][3]  ( .D(\in[3][3] ), .CK(clk), .Q(\add_in[3][3] ) );
  DFF_X1 \add_in_reg[3][2]  ( .D(\in[3][2] ), .CK(clk), .Q(\add_in[3][2] ) );
  DFF_X1 \add_in_reg[3][1]  ( .D(\in[3][1] ), .CK(clk), .Q(\add_in[3][1] ) );
  DFF_X1 \add_in_reg[3][0]  ( .D(\in[3][0] ), .CK(clk), .Q(\add_in[3][0] ) );
  DFF_X1 \add_in_reg[2][15]  ( .D(\in[2][15] ), .CK(clk), .Q(\add_in[2][15] )
         );
  DFF_X1 \add_in_reg[2][14]  ( .D(\in[2][14] ), .CK(clk), .Q(\add_in[2][14] )
         );
  DFF_X1 \add_in_reg[2][13]  ( .D(\in[2][13] ), .CK(clk), .Q(\add_in[2][13] )
         );
  DFF_X1 \add_in_reg[2][12]  ( .D(\in[2][12] ), .CK(clk), .Q(\add_in[2][12] )
         );
  DFF_X1 \add_in_reg[2][11]  ( .D(\in[2][11] ), .CK(clk), .Q(\add_in[2][11] )
         );
  DFF_X1 \add_in_reg[2][10]  ( .D(\in[2][10] ), .CK(clk), .Q(\add_in[2][10] )
         );
  DFF_X1 \add_in_reg[2][9]  ( .D(\in[2][9] ), .CK(clk), .Q(\add_in[2][9] ) );
  DFF_X1 \add_in_reg[2][8]  ( .D(\in[2][8] ), .CK(clk), .Q(\add_in[2][8] ) );
  DFF_X1 \add_in_reg[2][7]  ( .D(\in[2][7] ), .CK(clk), .Q(\add_in[2][7] ) );
  DFF_X1 \add_in_reg[2][6]  ( .D(\in[2][6] ), .CK(clk), .Q(\add_in[2][6] ) );
  DFF_X1 \add_in_reg[2][5]  ( .D(\in[2][5] ), .CK(clk), .Q(\add_in[2][5] ) );
  DFF_X1 \add_in_reg[2][4]  ( .D(\in[2][4] ), .CK(clk), .Q(\add_in[2][4] ) );
  DFF_X1 \add_in_reg[2][3]  ( .D(\in[2][3] ), .CK(clk), .Q(\add_in[2][3] ) );
  DFF_X1 \add_in_reg[2][2]  ( .D(\in[2][2] ), .CK(clk), .Q(\add_in[2][2] ) );
  DFF_X1 \add_in_reg[2][1]  ( .D(\in[2][1] ), .CK(clk), .Q(\add_in[2][1] ) );
  DFF_X1 \add_in_reg[2][0]  ( .D(\in[2][0] ), .CK(clk), .Q(\add_in[2][0] ) );
  DFF_X1 \add_in_reg[1][15]  ( .D(\in[1][15] ), .CK(clk), .Q(\add_in[1][15] )
         );
  DFF_X1 \add_in_reg[1][14]  ( .D(\in[1][14] ), .CK(clk), .Q(\add_in[1][14] )
         );
  DFF_X1 \add_in_reg[1][13]  ( .D(\in[1][13] ), .CK(clk), .Q(\add_in[1][13] )
         );
  DFF_X1 \add_in_reg[1][12]  ( .D(\in[1][12] ), .CK(clk), .Q(\add_in[1][12] )
         );
  DFF_X1 \add_in_reg[1][11]  ( .D(\in[1][11] ), .CK(clk), .Q(\add_in[1][11] )
         );
  DFF_X1 \add_in_reg[1][10]  ( .D(\in[1][10] ), .CK(clk), .Q(\add_in[1][10] )
         );
  DFF_X1 \add_in_reg[1][9]  ( .D(\in[1][9] ), .CK(clk), .Q(\add_in[1][9] ) );
  DFF_X1 \add_in_reg[1][8]  ( .D(\in[1][8] ), .CK(clk), .Q(\add_in[1][8] ) );
  DFF_X1 \add_in_reg[1][7]  ( .D(\in[1][7] ), .CK(clk), .Q(\add_in[1][7] ) );
  DFF_X1 \add_in_reg[1][6]  ( .D(\in[1][6] ), .CK(clk), .Q(\add_in[1][6] ) );
  DFF_X1 \add_in_reg[1][5]  ( .D(\in[1][5] ), .CK(clk), .Q(\add_in[1][5] ) );
  DFF_X1 \add_in_reg[1][4]  ( .D(\in[1][4] ), .CK(clk), .Q(\add_in[1][4] ) );
  DFF_X1 \add_in_reg[1][3]  ( .D(\in[1][3] ), .CK(clk), .Q(\add_in[1][3] ) );
  DFF_X1 \add_in_reg[1][2]  ( .D(\in[1][2] ), .CK(clk), .Q(\add_in[1][2] ) );
  DFF_X1 \add_in_reg[1][1]  ( .D(\in[1][1] ), .CK(clk), .Q(\add_in[1][1] ) );
  DFF_X1 \add_in_reg[1][0]  ( .D(\in[1][0] ), .CK(clk), .Q(\add_in[1][0] ) );
  DFF_X1 \add_in_reg[0][15]  ( .D(\in[0][15] ), .CK(clk), .Q(\add_in[0][15] )
         );
  DFF_X1 \add_in_reg[0][11]  ( .D(\in[0][11] ), .CK(clk), .Q(\add_in[0][11] )
         );
  DFF_X1 \add_in_reg[0][10]  ( .D(\in[0][10] ), .CK(clk), .Q(\add_in[0][10] )
         );
  DFF_X1 \add_in_reg[0][9]  ( .D(\in[0][9] ), .CK(clk), .Q(\add_in[0][9] ) );
  DFF_X1 \add_in_reg[0][8]  ( .D(\in[0][8] ), .CK(clk), .Q(\add_in[0][8] ) );
  DFF_X1 \add_in_reg[0][7]  ( .D(\in[0][7] ), .CK(clk), .Q(\add_in[0][7] ) );
  DFF_X1 \add_in_reg[0][6]  ( .D(\in[0][6] ), .CK(clk), .Q(\add_in[0][6] ) );
  DFF_X1 \add_in_reg[0][5]  ( .D(\in[0][5] ), .CK(clk), .Q(\add_in[0][5] ) );
  DFF_X1 \add_in_reg[0][4]  ( .D(\in[0][4] ), .CK(clk), .Q(\add_in[0][4] ) );
  DFF_X1 \add_in_reg[0][3]  ( .D(\in[0][3] ), .CK(clk), .Q(\add_in[0][3] ) );
  DFF_X1 \add_in_reg[0][2]  ( .D(\in[0][2] ), .CK(clk), .Q(\add_in[0][2] ) );
  DFF_X1 \add_in_reg[0][1]  ( .D(\in[0][1] ), .CK(clk), .Q(\add_in[0][1] ) );
  DFF_X1 \add_in_reg[0][0]  ( .D(\in[0][0] ), .CK(clk), .Q(\add_in[0][0] ) );
  add_layer_WIDTH16_6 \genblk2.genblk1[0].add_two_number  ( .clk(clk), .a({
        \add_in[0][15] , \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , 
        \add_in[0][11] , \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , 
        \add_in[0][7] , \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , 
        \add_in[0][3] , \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .b({
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), 
        .out({\genblk2.inter[0][15] , \genblk2.inter[0][14] , 
        \genblk2.inter[0][13] , \genblk2.inter[0][12] , \genblk2.inter[0][11] , 
        \genblk2.inter[0][10] , \genblk2.inter[0][9] , \genblk2.inter[0][8] , 
        \genblk2.inter[0][7] , \genblk2.inter[0][6] , \genblk2.inter[0][5] , 
        \genblk2.inter[0][4] , \genblk2.inter[0][3] , \genblk2.inter[0][2] , 
        \genblk2.inter[0][1] , \genblk2.inter[0][0] }) );
  add_layer_WIDTH16_5 \genblk2.genblk1[1].add_two_number  ( .clk(clk), .a({
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .b({
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), 
        .out({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE2_WIDTH16_1 \genblk2.next_layer  ( .clk(clk), 
        .in({\genblk2.inter[1][15] , \genblk2.inter[1][14] , 
        \genblk2.inter[1][13] , \genblk2.inter[1][12] , \genblk2.inter[1][11] , 
        \genblk2.inter[1][10] , \genblk2.inter[1][9] , \genblk2.inter[1][8] , 
        \genblk2.inter[1][7] , \genblk2.inter[1][6] , \genblk2.inter[1][5] , 
        \genblk2.inter[1][4] , \genblk2.inter[1][3] , \genblk2.inter[1][2] , 
        \genblk2.inter[1][1] , \genblk2.inter[1][0] , \genblk2.inter[0][15] , 
        \genblk2.inter[0][14] , \genblk2.inter[0][13] , \genblk2.inter[0][12] , 
        \genblk2.inter[0][11] , \genblk2.inter[0][10] , \genblk2.inter[0][9] , 
        \genblk2.inter[0][8] , \genblk2.inter[0][7] , \genblk2.inter[0][6] , 
        \genblk2.inter[0][5] , \genblk2.inter[0][4] , \genblk2.inter[0][3] , 
        \genblk2.inter[0][2] , \genblk2.inter[0][1] , \genblk2.inter[0][0] }), 
        .out(out) );
  DFF_X1 \add_in_reg[0][14]  ( .D(\in[0][14] ), .CK(clk), .Q(\add_in[0][14] )
         );
  DFF_X1 \add_in_reg[0][13]  ( .D(\in[0][13] ), .CK(clk), .Q(\add_in[0][13] )
         );
  DFF_X1 \add_in_reg[0][12]  ( .D(\in[0][12] ), .CK(clk), .Q(\add_in[0][12] )
         );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_1 ( clk, 
    .a({\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , 
        \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , 
        \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , 
        \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input clk, \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] ,
         \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] ,
         \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] ,
         \mult_out[3][6] , \mult_out[3][5] , \mult_out[3][4] ,
         \mult_out[3][3] , \mult_out[3][2] , \mult_out[3][1] ,
         \mult_out[3][0] , \mult_out[2][15] , \mult_out[2][14] ,
         \mult_out[2][13] , \mult_out[2][12] , \mult_out[2][11] ,
         \mult_out[2][10] , \mult_out[2][9] , \mult_out[2][8] ,
         \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] ,
         \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] ,
         \mult_out[2][1] , \mult_out[2][0] , \mult_out[1][15] ,
         \mult_out[1][14] , \mult_out[1][13] , \mult_out[1][12] ,
         \mult_out[1][11] , \mult_out[1][10] , \mult_out[1][9] ,
         \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] ,
         \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] ,
         \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] ,
         \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] ,
         \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] ,
         \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] ,
         \mult_out[0][6] , \mult_out[0][5] , \mult_out[0][4] ,
         \mult_out[0][3] , \mult_out[0][2] , \mult_out[0][1] ,
         \mult_out[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4 \genblk1[0].mult  ( .clk(clk), .ia(
        {\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , 
        \a[0][1] , \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , 
        \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3 \genblk1[1].mult  ( .clk(clk), .ia(
        {\a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , 
        \a[1][1] , \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({
        \mult_out[1][15] , \mult_out[1][14] , \mult_out[1][13] , 
        \mult_out[1][12] , \mult_out[1][11] , \mult_out[1][10] , 
        \mult_out[1][9] , \mult_out[1][8] , \mult_out[1][7] , \mult_out[1][6] , 
        \mult_out[1][5] , \mult_out[1][4] , \mult_out[1][3] , \mult_out[1][2] , 
        \mult_out[1][1] , \mult_out[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2 \genblk1[2].mult  ( .clk(clk), .ia(
        {\a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , 
        \a[2][1] , \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({
        \mult_out[2][15] , \mult_out[2][14] , \mult_out[2][13] , 
        \mult_out[2][12] , \mult_out[2][11] , \mult_out[2][10] , 
        \mult_out[2][9] , \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , 
        \mult_out[2][5] , \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , 
        \mult_out[2][1] , \mult_out[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1 \genblk1[3].mult  ( .clk(clk), .ia(
        {\a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , 
        \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_INTERREG1_1 add ( .clk(clk), .in({
        \mult_out[3][15] , \mult_out[3][14] , \mult_out[3][13] , 
        \mult_out[3][12] , \mult_out[3][11] , \mult_out[3][10] , 
        \mult_out[3][9] , \mult_out[3][8] , \mult_out[3][7] , \mult_out[3][6] , 
        \mult_out[3][5] , \mult_out[3][4] , \mult_out[3][3] , \mult_out[3][2] , 
        \mult_out[3][1] , \mult_out[3][0] , \mult_out[2][15] , 
        \mult_out[2][14] , \mult_out[2][13] , \mult_out[2][12] , 
        \mult_out[2][11] , \mult_out[2][10] , \mult_out[2][9] , 
        \mult_out[2][8] , \mult_out[2][7] , \mult_out[2][6] , \mult_out[2][5] , 
        \mult_out[2][4] , \mult_out[2][3] , \mult_out[2][2] , \mult_out[2][1] , 
        \mult_out[2][0] , \mult_out[1][15] , \mult_out[1][14] , 
        \mult_out[1][13] , \mult_out[1][12] , \mult_out[1][11] , 
        \mult_out[1][10] , \mult_out[1][9] , \mult_out[1][8] , 
        \mult_out[1][7] , \mult_out[1][6] , \mult_out[1][5] , \mult_out[1][4] , 
        \mult_out[1][3] , \mult_out[1][2] , \mult_out[1][1] , \mult_out[1][0] , 
        \mult_out[0][15] , \mult_out[0][14] , \mult_out[0][13] , 
        \mult_out[0][12] , \mult_out[0][11] , \mult_out[0][10] , 
        \mult_out[0][9] , \mult_out[0][8] , \mult_out[0][7] , \mult_out[0][6] , 
        \mult_out[0][5] , \mult_out[0][4] , \mult_out[0][3] , \mult_out[0][2] , 
        \mult_out[0][1] , \mult_out[0][0] }), .out(y) );
endmodule


module data_path_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_DELAY2 ( clk, 
        en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay, of_a, 
        of_x, of_y, of_delay, data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay;
  output of_a, of_x, of_y, of_delay;
  wire   N24, N25, \a[15][7] , \a[15][6] , \a[15][5] , \a[15][4] , \a[15][3] ,
         \a[15][2] , \a[15][1] , \a[15][0] , \a[14][7] , \a[14][6] ,
         \a[14][5] , \a[14][4] , \a[14][3] , \a[14][2] , \a[14][1] ,
         \a[14][0] , \a[13][7] , \a[13][6] , \a[13][5] , \a[13][4] ,
         \a[13][3] , \a[13][2] , \a[13][1] , \a[13][0] , \a[12][7] ,
         \a[12][6] , \a[12][5] , \a[12][4] , \a[12][3] , \a[12][2] ,
         \a[12][1] , \a[12][0] , \a[11][7] , \a[11][6] , \a[11][5] ,
         \a[11][4] , \a[11][3] , \a[11][2] , \a[11][1] , \a[11][0] ,
         \a[10][7] , \a[10][6] , \a[10][5] , \a[10][4] , \a[10][3] ,
         \a[10][2] , \a[10][1] , \a[10][0] , \a[9][7] , \a[9][6] , \a[9][5] ,
         \a[9][4] , \a[9][3] , \a[9][2] , \a[9][1] , \a[9][0] , \a[8][7] ,
         \a[8][6] , \a[8][5] , \a[8][4] , \a[8][3] , \a[8][2] , \a[8][1] ,
         \a[8][0] , \a[7][7] , \a[7][6] , \a[7][5] , \a[7][4] , \a[7][3] ,
         \a[7][2] , \a[7][1] , \a[7][0] , \a[6][7] , \a[6][6] , \a[6][5] ,
         \a[6][4] , \a[6][3] , \a[6][2] , \a[6][1] , \a[6][0] , \a[5][7] ,
         \a[5][6] , \a[5][5] , \a[5][4] , \a[5][3] , \a[5][2] , \a[5][1] ,
         \a[5][0] , \a[4][7] , \a[4][6] , \a[4][5] , \a[4][4] , \a[4][3] ,
         \a[4][2] , \a[4][1] , \a[4][0] , \a[3][7] , \a[3][6] , \a[3][5] ,
         \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , \a[3][0] , \a[2][7] ,
         \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , \a[2][1] ,
         \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] ,
         \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , \a[0][6] , \a[0][5] ,
         \a[0][4] , \a[0][2] , \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] ,
         \x[3][5] , \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] ,
         \x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] ,
         \x[2][1] , \x[2][0] , \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] ,
         \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] ,
         \x[0][5] , \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ,
         \y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] , \y[3][11] ,
         \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] , \y[3][5] ,
         \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] , \y[2][15] ,
         \y[2][14] , \y[2][13] , \y[2][12] , \y[2][11] , \y[2][10] , \y[2][9] ,
         \y[2][8] , \y[2][7] , \y[2][6] , \y[2][5] , \y[2][4] , \y[2][3] ,
         \y[2][2] , \y[2][1] , \y[2][0] , \y[1][15] , \y[1][14] , \y[1][13] ,
         \y[1][12] , \y[1][11] , \y[1][10] , \y[1][9] , \y[1][8] , \y[1][7] ,
         \y[1][6] , \y[1][5] , \y[1][4] , \y[1][3] , \y[1][2] , \y[1][1] ,
         \y[1][0] , \y[0][15] , \y[0][14] , \y[0][13] , \y[0][12] , \y[0][11] ,
         \y[0][10] , \y[0][9] , \y[0][8] , \y[0][7] , \y[0][6] , \y[0][5] ,
         \y[0][4] , \y[0][3] , \y[0][2] , \y[0][1] , \y[0][0] , N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N89,
         N91, N92, N96, N97, N101, N102, N108, N109, N110, N114, N115, N116,
         n9, n10, n12, n15, n16, n19, n20, n21, n32, n33, n41, n42, n43, n44,
         n52, n53, n54, n62, n63, n64, n72, n73, n74, n82, n83, n91, n92, n100,
         n101, n102, n110, n111, n119, n120, n128, n129, n137, n138, n146,
         n147, n155, n156, n157, n165, n166, n174, n175, n176, n184, n185,
         n186, n194, n195, n203, n204, n212, n213, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n1, n2, n3, n4, n5, n6, n7,
         n8, n11, n13, n14, n17, n18, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n34, n35, n36, n37, n38, n39, n40, n45, n46, n47, n48, n49,
         n50, n51, n55, n56, n57, n58, n59, n60, n61, n65, n66, n67, n68, n69,
         n70, n71, n75, n76, n77, n78, n79, n80, n81, n84, n85, n86, n87, n88,
         n89, n90, n93, n94, n95, n96, n97, n98, n99, n103, n104, n105, n106,
         n107, n108, n109, n112, n113, n114, n115, n116, n117, n118, n121,
         n122, n123, n124, n125, n126, n127, n130, n131, n132, n133, n134,
         n135, n136, n139, n140, n141, n142, n143, n144, n145, n148, n149,
         n150, n151, n152, n153, n154, n158, n159, n160, n161, n162, n163,
         n164, n167, n168, n169, n170, n171, n172, n173, n177, n178, n179,
         n180, n181, n182, n183, n187, n188, n189, n190, n191, n192, n193,
         n196, n197, n198, n199, n200, n201, n202, n205, n206, n207, n208,
         n209, n210, n211, n214, n215, n216, n217, n218, n219, n220, n230,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444;
  wire   [3:0] addr_a;
  wire   [1:0] addr_x;
  wire   [3:0] delay_timer;
  assign of_a = N114;
  assign of_x = N115;
  assign of_y = N116;

  DFF_X1 \data_out_reg[15]  ( .D(N68), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N69), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N70), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N71), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N72), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N73), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N74), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N75), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N76), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N77), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N78), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N79), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N80), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N81), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N82), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N83), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \addr_a_reg[0]  ( .D(N89), .CK(clk), .Q(addr_a[0]) );
  DFF_X1 \addr_a_reg[1]  ( .D(n440), .CK(clk), .Q(addr_a[1]), .QN(n12) );
  DFF_X1 \addr_a_reg[2]  ( .D(N91), .CK(clk), .Q(addr_a[2]), .QN(n10) );
  DFF_X1 \addr_a_reg[3]  ( .D(N92), .CK(clk), .Q(addr_a[3]), .QN(n9) );
  DFF_X1 \a_reg[3][6]  ( .D(n356), .CK(clk), .Q(\a[3][6] ) );
  DFF_X1 \a_reg[3][4]  ( .D(n358), .CK(clk), .Q(\a[3][4] ) );
  DFF_X1 \a_reg[3][2]  ( .D(n360), .CK(clk), .Q(\a[3][2] ) );
  DFF_X1 \a_reg[3][0]  ( .D(n362), .CK(clk), .Q(\a[3][0] ) );
  DFF_X1 \a_reg[2][6]  ( .D(n364), .CK(clk), .Q(\a[2][6] ) );
  DFF_X1 \a_reg[2][4]  ( .D(n366), .CK(clk), .Q(\a[2][4] ) );
  DFF_X1 \a_reg[2][2]  ( .D(n368), .CK(clk), .Q(\a[2][2] ) );
  DFF_X1 \a_reg[2][0]  ( .D(n370), .CK(clk), .Q(\a[2][0] ) );
  DFF_X1 \a_reg[1][6]  ( .D(n372), .CK(clk), .Q(\a[1][6] ), .QN(n117) );
  DFF_X1 \a_reg[1][4]  ( .D(n374), .CK(clk), .Q(\a[1][4] ) );
  DFF_X1 \a_reg[1][2]  ( .D(n376), .CK(clk), .Q(\a[1][2] ) );
  DFF_X1 \a_reg[1][0]  ( .D(n378), .CK(clk), .Q(\a[1][0] ) );
  DFF_X1 \a_reg[0][6]  ( .D(n380), .CK(clk), .Q(\a[0][6] ) );
  DFF_X1 \a_reg[0][4]  ( .D(n382), .CK(clk), .Q(\a[0][4] ), .QN(n14) );
  DFF_X1 \a_reg[0][2]  ( .D(n384), .CK(clk), .Q(\a[0][2] ) );
  DFF_X1 \a_reg[0][0]  ( .D(n386), .CK(clk), .Q(\a[0][0] ) );
  DFF_X1 \a_reg[11][7]  ( .D(n291), .CK(clk), .Q(\a[11][7] ) );
  DFF_X1 \a_reg[11][6]  ( .D(n292), .CK(clk), .Q(\a[11][6] ) );
  DFF_X1 \a_reg[11][4]  ( .D(n294), .CK(clk), .Q(\a[11][4] ) );
  DFF_X1 \a_reg[11][3]  ( .D(n295), .CK(clk), .Q(\a[11][3] ), .QN(n105) );
  DFF_X1 \a_reg[11][2]  ( .D(n296), .CK(clk), .Q(\a[11][2] ) );
  DFF_X1 \a_reg[11][0]  ( .D(n298), .CK(clk), .Q(\a[11][0] ) );
  DFF_X1 \a_reg[10][6]  ( .D(n300), .CK(clk), .Q(\a[10][6] ) );
  DFF_X1 \a_reg[10][4]  ( .D(n302), .CK(clk), .Q(\a[10][4] ) );
  DFF_X1 \a_reg[10][2]  ( .D(n304), .CK(clk), .Q(\a[10][2] ) );
  DFF_X1 \a_reg[10][1]  ( .D(n305), .CK(clk), .Q(\a[10][1] ), .QN(n31) );
  DFF_X1 \a_reg[10][0]  ( .D(n306), .CK(clk), .Q(\a[10][0] ) );
  DFF_X1 \a_reg[9][6]  ( .D(n308), .CK(clk), .Q(\a[9][6] ), .QN(n78) );
  DFF_X1 \a_reg[9][4]  ( .D(n310), .CK(clk), .Q(\a[9][4] ) );
  DFF_X1 \a_reg[9][2]  ( .D(n312), .CK(clk), .Q(\a[9][2] ) );
  DFF_X1 \a_reg[9][0]  ( .D(n314), .CK(clk), .Q(\a[9][0] ) );
  DFF_X1 \a_reg[8][6]  ( .D(n316), .CK(clk), .Q(\a[8][6] ), .QN(n27) );
  DFF_X1 \a_reg[8][4]  ( .D(n318), .CK(clk), .Q(\a[8][4] ) );
  DFF_X1 \a_reg[8][3]  ( .D(n319), .CK(clk), .Q(\a[8][3] ), .QN(n29) );
  DFF_X1 \a_reg[8][2]  ( .D(n320), .CK(clk), .Q(\a[8][2] ), .QN(n49) );
  DFF_X1 \a_reg[8][0]  ( .D(n322), .CK(clk), .Q(\a[8][0] ) );
  DFF_X1 \a_reg[14][6]  ( .D(n268), .CK(clk), .Q(\a[14][6] ) );
  DFF_X1 \a_reg[14][4]  ( .D(n270), .CK(clk), .Q(\a[14][4] ) );
  DFF_X1 \a_reg[14][2]  ( .D(n272), .CK(clk), .Q(\a[14][2] ), .QN(n11) );
  DFF_X1 \a_reg[14][0]  ( .D(n274), .CK(clk), .Q(\a[14][0] ) );
  DFF_X1 \a_reg[13][7]  ( .D(n275), .CK(clk), .Q(\a[13][7] ), .QN(n67) );
  DFF_X1 \a_reg[13][6]  ( .D(n276), .CK(clk), .Q(\a[13][6] ) );
  DFF_X1 \a_reg[13][4]  ( .D(n278), .CK(clk), .Q(\a[13][4] ) );
  DFF_X1 \a_reg[13][2]  ( .D(n280), .CK(clk), .Q(\a[13][2] ) );
  DFF_X1 \a_reg[13][0]  ( .D(n282), .CK(clk), .Q(\a[13][0] ) );
  DFF_X1 \a_reg[12][5]  ( .D(n285), .CK(clk), .Q(\a[12][5] ), .QN(n403) );
  DFF_X1 \a_reg[12][4]  ( .D(n286), .CK(clk), .Q(\a[12][4] ) );
  DFF_X1 \a_reg[12][2]  ( .D(n288), .CK(clk), .Q(\a[12][2] ) );
  DFF_X1 \a_reg[12][0]  ( .D(n290), .CK(clk), .Q(\a[12][0] ) );
  DFF_X1 \a_reg[6][6]  ( .D(n332), .CK(clk), .Q(\a[6][6] ) );
  DFF_X1 \a_reg[6][4]  ( .D(n334), .CK(clk), .Q(\a[6][4] ) );
  DFF_X1 \a_reg[6][2]  ( .D(n336), .CK(clk), .Q(\a[6][2] ) );
  DFF_X1 \a_reg[6][0]  ( .D(n338), .CK(clk), .Q(\a[6][0] ) );
  DFF_X1 \a_reg[5][7]  ( .D(n339), .CK(clk), .Q(\a[5][7] ) );
  DFF_X1 \a_reg[5][6]  ( .D(n340), .CK(clk), .Q(\a[5][6] ) );
  DFF_X1 \a_reg[5][4]  ( .D(n342), .CK(clk), .Q(\a[5][4] ) );
  DFF_X1 \a_reg[5][2]  ( .D(n344), .CK(clk), .Q(\a[5][2] ) );
  DFF_X1 \a_reg[5][0]  ( .D(n346), .CK(clk), .Q(\a[5][0] ) );
  DFF_X1 \a_reg[4][6]  ( .D(n348), .CK(clk), .Q(\a[4][6] ) );
  DFF_X1 \a_reg[4][4]  ( .D(n350), .CK(clk), .Q(\a[4][4] ) );
  DFF_X1 \a_reg[4][2]  ( .D(n352), .CK(clk), .Q(\a[4][2] ), .QN(n18) );
  DFF_X1 \a_reg[4][0]  ( .D(n354), .CK(clk), .Q(\a[4][0] ) );
  DFF_X1 \a_reg[7][7]  ( .D(n323), .CK(clk), .Q(\a[7][7] ) );
  DFF_X1 \a_reg[7][6]  ( .D(n324), .CK(clk), .Q(\a[7][6] ) );
  DFF_X1 \a_reg[7][4]  ( .D(n326), .CK(clk), .Q(\a[7][4] ) );
  DFF_X1 \a_reg[7][2]  ( .D(n328), .CK(clk), .Q(\a[7][2] ) );
  DFF_X1 \a_reg[7][0]  ( .D(n330), .CK(clk), .Q(\a[7][0] ) );
  DFF_X1 \a_reg[15][6]  ( .D(n260), .CK(clk), .Q(\a[15][6] ) );
  DFF_X1 \a_reg[15][4]  ( .D(n262), .CK(clk), .Q(\a[15][4] ) );
  DFF_X1 \a_reg[15][2]  ( .D(n264), .CK(clk), .Q(\a[15][2] ) );
  DFF_X1 \a_reg[15][0]  ( .D(n266), .CK(clk), .Q(\a[15][0] ) );
  DFF_X1 \addr_x_reg[0]  ( .D(N96), .CK(clk), .Q(addr_x[0]), .QN(n16) );
  DFF_X1 \addr_x_reg[1]  ( .D(N97), .CK(clk), .Q(addr_x[1]), .QN(n15) );
  DFF_X1 \x_reg[2][6]  ( .D(n236), .CK(clk), .Q(\x[2][6] ), .QN(n39) );
  DFF_X1 \x_reg[2][5]  ( .D(n237), .CK(clk), .Q(\x[2][5] ), .QN(n47) );
  DFF_X1 \x_reg[2][4]  ( .D(n238), .CK(clk), .Q(\x[2][4] ) );
  DFF_X1 \x_reg[2][2]  ( .D(n240), .CK(clk), .Q(\x[2][2] ) );
  DFF_X1 \x_reg[2][0]  ( .D(n242), .CK(clk), .Q(\x[2][0] ), .QN(n35) );
  DFF_X1 \x_reg[0][4]  ( .D(n254), .CK(clk), .Q(\x[0][4] ), .QN(n125) );
  DFF_X1 \x_reg[0][2]  ( .D(n256), .CK(clk), .Q(\x[0][2] ), .QN(n86) );
  DFF_X1 \x_reg[0][0]  ( .D(n258), .CK(clk), .Q(\x[0][0] ) );
  DFF_X1 \x_reg[1][7]  ( .D(n243), .CK(clk), .Q(\x[1][7] ), .QN(n121) );
  DFF_X1 \x_reg[1][0]  ( .D(n250), .CK(clk), .Q(\x[1][0] ), .QN(n23) );
  DFF_X1 \x_reg[3][7]  ( .D(n431), .CK(clk), .Q(\x[3][7] ), .QN(n80) );
  DFF_X1 \x_reg[3][2]  ( .D(n436), .CK(clk), .Q(\x[3][2] ), .QN(n96) );
  DFF_X1 \x_reg[3][0]  ( .D(n438), .CK(clk), .Q(\x[3][0] ) );
  DFF_X1 \addr_y_reg[1]  ( .D(N102), .CK(clk), .Q(N25), .QN(n4) );
  DFF_X1 \delay_timer_reg[0]  ( .D(N108), .CK(clk), .Q(delay_timer[0]), .QN(
        n21) );
  DFF_X1 \delay_timer_reg[1]  ( .D(N109), .CK(clk), .Q(delay_timer[1]), .QN(
        n20) );
  DFF_X1 \delay_timer_reg[2]  ( .D(N110), .CK(clk), .Q(delay_timer[2]), .QN(
        n19) );
  DFF_X1 \delay_timer_reg[3]  ( .D(n442), .CK(clk), .Q(delay_timer[3]) );
  NAND3_X1 U394 ( .A1(delay_timer[0]), .A2(n443), .A3(delay_timer[1]), .ZN(
        n231) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_0 \genblk1[0].element  ( 
        .clk(clk), .a({n154, \a[3][6] , n406, \a[3][4] , n114, \a[3][2] , 
        \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , 
        \a[2][3] , \a[2][2] , n230, \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , 
        \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , 
        \a[0][6] , n95, \a[0][4] , n408, \a[0][2] , \a[0][1] , \a[0][0] }), 
        .x({n81, \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , n97, \x[3][1] , 
        \x[3][0] , n116, n40, n48, n214, n89, n215, n159, n36, \x[1][7] , n75, 
        \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] , n124, 
        n85, n61, n126, \x[0][3] , n87, \x[0][1] , \x[0][0] }), .y({\y[0][15] , 
        \y[0][14] , \y[0][13] , \y[0][12] , \y[0][11] , \y[0][10] , \y[0][9] , 
        \y[0][8] , \y[0][7] , \y[0][6] , \y[0][5] , \y[0][4] , \y[0][3] , 
        \y[0][2] , \y[0][1] , \y[0][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_3 \genblk1[1].element  ( 
        .clk(clk), .a({\a[7][7] , \a[7][6] , \a[7][5] , \a[7][4] , n390, 
        \a[7][2] , n152, \a[7][0] , \a[6][7] , \a[6][6] , n394, \a[6][4] , 
        \a[6][3] , \a[6][2] , \a[6][1] , \a[6][0] , \a[5][7] , \a[5][6] , n402, 
        \a[5][4] , \a[5][3] , \a[5][2] , \a[5][1] , \a[5][0] , n108, \a[4][6] , 
        \a[4][5] , \a[4][4] , \a[4][3] , \a[4][2] , \a[4][1] , \a[4][0] }), 
        .x({\x[3][7] , n70, \x[3][5] , \x[3][4] , n55, n97, n217, \x[3][0] , 
        n116, n40, n48, n214, n89, n215, \x[2][1] , \x[2][0] , n122, \x[1][6] , 
        \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , n130, n24, \x[0][7] , 
        \x[0][6] , \x[0][5] , n126, \x[0][3] , n87, n400, \x[0][0] }), .y({
        \y[1][15] , \y[1][14] , \y[1][13] , \y[1][12] , \y[1][11] , \y[1][10] , 
        \y[1][9] , \y[1][8] , \y[1][7] , \y[1][6] , \y[1][5] , \y[1][4] , 
        \y[1][3] , \y[1][2] , \y[1][1] , \y[1][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_2 \genblk1[2].element  ( 
        .clk(clk), .a({\a[11][7] , \a[11][6] , n136, \a[11][4] , \a[11][3] , 
        \a[11][2] , \a[11][1] , \a[11][0] , \a[10][7] , \a[10][6] , n148, 
        \a[10][4] , \a[10][3] , \a[10][2] , \a[10][1] , \a[10][0] , \a[9][7] , 
        \a[9][6] , n142, \a[9][4] , \a[9][3] , \a[9][2] , \a[9][1] , \a[9][0] , 
        \a[8][7] , \a[8][6] , n388, \a[8][4] , \a[8][3] , \a[8][2] , \a[8][1] , 
        \a[8][0] }), .x({n81, n70, \x[3][5] , \x[3][4] , n55, \x[3][2] , 
        \x[3][1] , \x[3][0] , \x[2][7] , n40, n48, n214, \x[2][3] , n215, n159, 
        \x[2][0] , \x[1][7] , n75, n59, n38, \x[1][3] , n66, \x[1][1] , 
        \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , 
        \x[0][2] , \x[0][1] , \x[0][0] }), .y({\y[2][15] , \y[2][14] , 
        \y[2][13] , \y[2][12] , \y[2][11] , \y[2][10] , \y[2][9] , \y[2][8] , 
        \y[2][7] , \y[2][6] , \y[2][5] , \y[2][4] , \y[2][3] , \y[2][2] , 
        \y[2][1] , \y[2][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_1 \genblk1[3].element  ( 
        .clk(clk), .a({n26, \a[15][6] , \a[15][5] , \a[15][4] , \a[15][3] , 
        \a[15][2] , \a[15][1] , \a[15][0] , n46, \a[14][6] , \a[14][5] , 
        \a[14][4] , \a[14][3] , \a[14][2] , \a[14][1] , \a[14][0] , n68, 
        \a[13][6] , \a[13][5] , \a[13][4] , n140, \a[13][2] , \a[13][1] , 
        \a[13][0] , n167, \a[12][6] , n404, \a[12][4] , \a[12][3] , \a[12][2] , 
        n163, \a[12][0] }), .x({n81, \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , n214, n89, n215, n159, \x[2][0] , n122, n75, n59, n38, n396, 
        n66, n130, \x[1][0] , n124, n85, n61, \x[0][4] , \x[0][3] , n87, 
        \x[0][1] , \x[0][0] }), .y({\y[3][15] , \y[3][14] , \y[3][13] , 
        \y[3][12] , \y[3][11] , \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , 
        \y[3][6] , \y[3][5] , \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , 
        \y[3][0] }) );
  DFF_X2 \x_reg[1][1]  ( .D(n249), .CK(clk), .Q(\x[1][1] ), .QN(n127) );
  DFF_X2 \x_reg[0][3]  ( .D(n255), .CK(clk), .Q(\x[0][3] ) );
  DFF_X1 \a_reg[0][3]  ( .D(n383), .CK(clk), .QN(n407) );
  DFF_X1 \a_reg[3][5]  ( .D(n357), .CK(clk), .Q(\a[3][5] ), .QN(n405) );
  DFF_X1 \a_reg[8][1]  ( .D(n321), .CK(clk), .Q(\a[8][1] ), .QN(n103) );
  DFF_X1 \a_reg[5][1]  ( .D(n345), .CK(clk), .Q(\a[5][1] ) );
  DFF_X1 \a_reg[5][5]  ( .D(n341), .CK(clk), .Q(\a[5][5] ), .QN(n401) );
  DFF_X1 \a_reg[9][1]  ( .D(n313), .CK(clk), .Q(\a[9][1] ), .QN(n90) );
  DFF_X2 \x_reg[0][1]  ( .D(n257), .CK(clk), .Q(\x[0][1] ), .QN(n399) );
  DFF_X1 \a_reg[15][1]  ( .D(n265), .CK(clk), .Q(\a[15][1] ) );
  DFF_X1 \a_reg[4][1]  ( .D(n353), .CK(clk), .Q(\a[4][1] ), .QN(n397) );
  DFF_X2 \x_reg[1][3]  ( .D(n247), .CK(clk), .Q(\x[1][3] ), .QN(n395) );
  DFF_X1 \a_reg[6][5]  ( .D(n333), .CK(clk), .Q(\a[6][5] ), .QN(n393) );
  DFF_X1 \a_reg[15][5]  ( .D(n261), .CK(clk), .Q(\a[15][5] ) );
  DFF_X1 \a_reg[2][5]  ( .D(n365), .CK(clk), .Q(\a[2][5] ) );
  DFF_X1 \a_reg[9][3]  ( .D(n311), .CK(clk), .Q(\a[9][3] ), .QN(n391) );
  DFF_X1 \a_reg[7][3]  ( .D(n327), .CK(clk), .Q(\a[7][3] ), .QN(n389) );
  DFF_X1 \a_reg[8][5]  ( .D(n317), .CK(clk), .Q(\a[8][5] ), .QN(n387) );
  DFF_X1 \a_reg[2][1]  ( .D(n369), .CK(clk), .Q(\a[2][1] ), .QN(n220) );
  DFF_X1 \a_reg[13][5]  ( .D(n277), .CK(clk), .Q(\a[13][5] ) );
  DFF_X2 \x_reg[3][4]  ( .D(n434), .CK(clk), .Q(\x[3][4] ) );
  DFF_X1 \a_reg[14][1]  ( .D(n273), .CK(clk), .Q(\a[14][1] ), .QN(n218) );
  DFF_X2 \x_reg[3][1]  ( .D(n437), .CK(clk), .Q(\x[3][1] ), .QN(n216) );
  DFF_X1 \a_reg[4][3]  ( .D(n351), .CK(clk), .Q(\a[4][3] ) );
  DFF_X1 \a_reg[12][3]  ( .D(n287), .CK(clk), .Q(\a[12][3] ), .QN(n7) );
  DFF_X1 \a_reg[13][1]  ( .D(n281), .CK(clk), .Q(\a[13][1] ) );
  DFF_X1 \a_reg[12][6]  ( .D(n284), .CK(clk), .Q(\a[12][6] ) );
  DFF_X1 \a_reg[12][7]  ( .D(n283), .CK(clk), .Q(\a[12][7] ), .QN(n164) );
  DFF_X2 \a_reg[10][3]  ( .D(n303), .CK(clk), .Q(\a[10][3] ) );
  DFF_X1 \a_reg[12][1]  ( .D(n289), .CK(clk), .Q(\a[12][1] ), .QN(n162) );
  DFF_X1 \a_reg[11][1]  ( .D(n297), .CK(clk), .Q(\a[11][1] ), .QN(n109) );
  DFF_X1 \a_reg[2][3]  ( .D(n367), .CK(clk), .Q(\a[2][3] ) );
  DFF_X1 \a_reg[7][5]  ( .D(n325), .CK(clk), .Q(\a[7][5] ), .QN(n160) );
  DFF_X1 \x_reg[2][1]  ( .D(n241), .CK(clk), .Q(\x[2][1] ), .QN(n158) );
  DFF_X1 \a_reg[14][3]  ( .D(n271), .CK(clk), .Q(\a[14][3] ) );
  DFF_X1 \a_reg[3][7]  ( .D(n355), .CK(clk), .Q(\a[3][7] ), .QN(n153) );
  DFF_X1 \a_reg[7][1]  ( .D(n329), .CK(clk), .Q(\a[7][1] ), .QN(n151) );
  DFF_X1 \a_reg[0][1]  ( .D(n385), .CK(clk), .Q(\a[0][1] ) );
  DFF_X1 \a_reg[10][5]  ( .D(n301), .CK(clk), .Q(\a[10][5] ), .QN(n145) );
  DFF_X1 \a_reg[9][5]  ( .D(n309), .CK(clk), .Q(\a[9][5] ), .QN(n141) );
  DFF_X1 \a_reg[13][3]  ( .D(n279), .CK(clk), .Q(\a[13][3] ), .QN(n139) );
  DFF_X1 \a_reg[14][5]  ( .D(n269), .CK(clk), .Q(\a[14][5] ) );
  DFF_X1 \a_reg[6][1]  ( .D(n337), .CK(clk), .Q(\a[6][1] ) );
  DFF_X1 \a_reg[11][5]  ( .D(n293), .CK(clk), .Q(\a[11][5] ), .QN(n135) );
  DFF_X1 \a_reg[1][7]  ( .D(n371), .CK(clk), .Q(\a[1][7] ) );
  DFF_X1 \a_reg[10][7]  ( .D(n299), .CK(clk), .Q(\a[10][7] ) );
  DFF_X1 \a_reg[5][3]  ( .D(n343), .CK(clk), .Q(\a[5][3] ), .QN(n133) );
  DFF_X1 \a_reg[9][7]  ( .D(n307), .CK(clk), .Q(\a[9][7] ), .QN(n131) );
  DFF_X1 \a_reg[6][3]  ( .D(n335), .CK(clk), .Q(\a[6][3] ) );
  DFF_X1 \a_reg[0][7]  ( .D(n379), .CK(clk), .Q(\a[0][7] ) );
  DFF_X1 \a_reg[1][1]  ( .D(n377), .CK(clk), .Q(\a[1][1] ), .QN(n409) );
  DFF_X1 \a_reg[3][1]  ( .D(n361), .CK(clk), .Q(\a[3][1] ), .QN(n76) );
  DFF_X1 \a_reg[1][5]  ( .D(n373), .CK(clk), .Q(\a[1][5] ), .QN(n56) );
  DFF_X2 \x_reg[3][5]  ( .D(n433), .CK(clk), .Q(\x[3][5] ) );
  DFF_X1 \x_reg[2][7]  ( .D(n235), .CK(clk), .Q(\x[2][7] ), .QN(n115) );
  DFF_X1 \a_reg[3][3]  ( .D(n359), .CK(clk), .Q(\a[3][3] ), .QN(n113) );
  DFF_X1 \a_reg[4][7]  ( .D(n347), .CK(clk), .Q(\a[4][7] ), .QN(n107) );
  DFF_X1 \a_reg[15][3]  ( .D(n263), .CK(clk), .Q(\a[15][3] ), .QN(n149) );
  DFF_X1 \a_reg[1][3]  ( .D(n375), .CK(clk), .Q(\a[1][3] ), .QN(n98) );
  DFF_X1 \a_reg[2][7]  ( .D(n363), .CK(clk), .Q(\a[2][7] ) );
  DFF_X1 \a_reg[8][7]  ( .D(n315), .CK(clk), .Q(\a[8][7] ) );
  DFF_X1 \a_reg[0][5]  ( .D(n381), .CK(clk), .Q(\a[0][5] ), .QN(n94) );
  DFF_X1 \x_reg[2][3]  ( .D(n239), .CK(clk), .Q(\x[2][3] ), .QN(n88) );
  DFF_X1 \x_reg[0][6]  ( .D(n252), .CK(clk), .Q(\x[0][6] ), .QN(n84) );
  DFF_X1 \x_reg[1][6]  ( .D(n244), .CK(clk), .Q(\x[1][6] ), .QN(n71) );
  DFF_X1 \x_reg[3][6]  ( .D(n432), .CK(clk), .Q(\x[3][6] ), .QN(n69) );
  DFF_X1 \x_reg[1][2]  ( .D(n248), .CK(clk), .Q(\x[1][2] ), .QN(n65) );
  DFF_X1 \x_reg[0][5]  ( .D(n253), .CK(clk), .Q(\x[0][5] ), .QN(n60) );
  DFF_X1 \x_reg[1][5]  ( .D(n245), .CK(clk), .Q(\x[1][5] ), .QN(n58) );
  DFF_X1 \x_reg[3][3]  ( .D(n435), .CK(clk), .Q(\x[3][3] ), .QN(n51) );
  DFF_X2 \x_reg[0][7]  ( .D(n251), .CK(clk), .Q(\x[0][7] ), .QN(n123) );
  DFF_X1 \a_reg[14][7]  ( .D(n267), .CK(clk), .Q(\a[14][7] ), .QN(n45) );
  DFF_X1 \x_reg[1][4]  ( .D(n246), .CK(clk), .Q(\x[1][4] ), .QN(n37) );
  DFF_X1 \a_reg[4][5]  ( .D(n349), .CK(clk), .Q(\a[4][5] ), .QN(n143) );
  DFF_X1 \a_reg[15][7]  ( .D(n259), .CK(clk), .Q(\a[15][7] ), .QN(n25) );
  DFF_X1 \addr_y_reg[0]  ( .D(N101), .CK(clk), .Q(N24), .QN(n210) );
  DFF_X2 \a_reg[6][7]  ( .D(n331), .CK(clk), .Q(\a[6][7] ) );
  INV_X2 U3 ( .A(n94), .ZN(n95) );
  INV_X2 U4 ( .A(n405), .ZN(n406) );
  INV_X1 U5 ( .A(n145), .ZN(n148) );
  INV_X1 U6 ( .A(n131), .ZN(n132) );
  INV_X1 U7 ( .A(n160), .ZN(n161) );
  AND2_X1 U8 ( .A1(N24), .A2(n4), .ZN(n1) );
  AND2_X1 U9 ( .A1(n4), .A2(n210), .ZN(n2) );
  AND2_X1 U10 ( .A1(N25), .A2(n210), .ZN(n3) );
  NOR3_X1 U11 ( .A1(n231), .A2(delay_timer[3]), .A3(n19), .ZN(n5) );
  CLKBUF_X1 U12 ( .A(n408), .Z(n6) );
  INV_X1 U13 ( .A(n7), .ZN(n8) );
  INV_X1 U14 ( .A(n11), .ZN(n13) );
  INV_X1 U15 ( .A(n14), .ZN(n17) );
  INV_X1 U16 ( .A(n18), .ZN(n22) );
  INV_X1 U17 ( .A(n23), .ZN(n24) );
  INV_X2 U18 ( .A(n25), .ZN(n26) );
  INV_X1 U19 ( .A(n27), .ZN(n28) );
  INV_X2 U20 ( .A(n121), .ZN(n122) );
  INV_X1 U21 ( .A(n29), .ZN(n30) );
  INV_X1 U22 ( .A(n31), .ZN(n34) );
  INV_X1 U23 ( .A(n35), .ZN(n36) );
  INV_X2 U24 ( .A(n37), .ZN(n38) );
  INV_X2 U25 ( .A(n39), .ZN(n40) );
  INV_X2 U26 ( .A(n45), .ZN(n46) );
  INV_X2 U27 ( .A(n47), .ZN(n48) );
  INV_X1 U28 ( .A(n49), .ZN(n50) );
  INV_X2 U29 ( .A(n51), .ZN(n55) );
  INV_X1 U30 ( .A(n56), .ZN(n57) );
  INV_X2 U31 ( .A(n58), .ZN(n59) );
  INV_X2 U32 ( .A(n60), .ZN(n61) );
  INV_X2 U33 ( .A(n65), .ZN(n66) );
  INV_X2 U34 ( .A(n67), .ZN(n68) );
  INV_X2 U35 ( .A(n69), .ZN(n70) );
  INV_X2 U36 ( .A(n71), .ZN(n75) );
  INV_X1 U37 ( .A(n76), .ZN(n77) );
  INV_X1 U38 ( .A(n78), .ZN(n79) );
  INV_X2 U39 ( .A(n80), .ZN(n81) );
  INV_X2 U40 ( .A(n84), .ZN(n85) );
  INV_X1 U41 ( .A(n133), .ZN(n134) );
  INV_X2 U42 ( .A(n86), .ZN(n87) );
  INV_X2 U43 ( .A(n88), .ZN(n89) );
  INV_X1 U44 ( .A(n90), .ZN(n93) );
  INV_X2 U45 ( .A(n96), .ZN(n97) );
  INV_X1 U46 ( .A(n98), .ZN(n99) );
  INV_X1 U47 ( .A(n103), .ZN(n104) );
  INV_X1 U48 ( .A(n105), .ZN(n106) );
  INV_X2 U49 ( .A(n107), .ZN(n108) );
  INV_X1 U50 ( .A(n109), .ZN(n112) );
  INV_X2 U51 ( .A(n113), .ZN(n114) );
  INV_X2 U52 ( .A(n115), .ZN(n116) );
  INV_X1 U53 ( .A(n117), .ZN(n118) );
  INV_X2 U54 ( .A(n123), .ZN(n124) );
  INV_X1 U55 ( .A(n391), .ZN(n392) );
  INV_X1 U56 ( .A(n397), .ZN(n398) );
  INV_X2 U57 ( .A(n125), .ZN(n126) );
  INV_X1 U58 ( .A(n218), .ZN(n219) );
  INV_X2 U59 ( .A(n127), .ZN(n130) );
  INV_X1 U60 ( .A(n162), .ZN(n163) );
  INV_X2 U61 ( .A(n135), .ZN(n136) );
  INV_X2 U62 ( .A(n139), .ZN(n140) );
  INV_X2 U63 ( .A(n141), .ZN(n142) );
  INV_X1 U64 ( .A(n143), .ZN(n144) );
  INV_X1 U65 ( .A(n149), .ZN(n150) );
  INV_X2 U66 ( .A(n151), .ZN(n152) );
  INV_X2 U67 ( .A(n153), .ZN(n154) );
  INV_X1 U68 ( .A(n220), .ZN(n230) );
  INV_X2 U69 ( .A(n158), .ZN(n159) );
  INV_X2 U70 ( .A(n164), .ZN(n167) );
  BUF_X4 U71 ( .A(\x[2][2] ), .Z(n215) );
  INV_X1 U72 ( .A(data_in[7]), .ZN(n444) );
  INV_X1 U73 ( .A(n210), .ZN(n211) );
  OAI21_X1 U74 ( .B1(n444), .B2(n119), .A(n120), .ZN(n243) );
  INV_X1 U75 ( .A(n227), .ZN(n440) );
  OAI21_X1 U76 ( .B1(n41), .B2(n52), .A(n441), .ZN(n227) );
  NOR4_X1 U77 ( .A1(delay_timer[3]), .A2(delay_timer[2]), .A3(delay_timer[1]), 
        .A4(n21), .ZN(of_delay) );
  NOR3_X1 U78 ( .A1(n225), .A2(n10), .A3(n9), .ZN(N114) );
  NOR2_X1 U79 ( .A1(n12), .A2(addr_a[0]), .ZN(n41) );
  AOI21_X1 U80 ( .B1(n20), .B2(n443), .A(N108), .ZN(n232) );
  AOI21_X1 U81 ( .B1(n441), .B2(n12), .A(N89), .ZN(n222) );
  NOR2_X1 U82 ( .A1(n15), .A2(n16), .ZN(N115) );
  NOR2_X1 U83 ( .A1(addr_a[0]), .A2(addr_a[1]), .ZN(n62) );
  OAI22_X1 U84 ( .A1(n232), .A2(n19), .B1(delay_timer[2]), .B2(n231), .ZN(N110) );
  OAI22_X1 U85 ( .A1(n222), .A2(n9), .B1(clr_addr_a), .B2(n223), .ZN(N92) );
  AOI22_X1 U86 ( .A1(n224), .A2(n430), .B1(addr_a[3]), .B2(n10), .ZN(n223) );
  NOR2_X1 U87 ( .A1(addr_a[3]), .A2(n10), .ZN(n224) );
  OAI22_X1 U88 ( .A1(n222), .A2(n10), .B1(n225), .B2(n226), .ZN(N91) );
  NAND2_X1 U89 ( .A1(n10), .A2(n441), .ZN(n226) );
  INV_X1 U90 ( .A(n228), .ZN(n442) );
  AOI21_X1 U91 ( .B1(n229), .B2(delay_timer[3]), .A(n5), .ZN(n228) );
  OAI21_X1 U92 ( .B1(clr_delay), .B2(delay_timer[2]), .A(n232), .ZN(n229) );
  OAI21_X1 U93 ( .B1(n444), .B2(n137), .A(n138), .ZN(n259) );
  OAI21_X1 U94 ( .B1(n444), .B2(n212), .A(n213), .ZN(n323) );
  OAI21_X1 U95 ( .B1(n444), .B2(n43), .A(n44), .ZN(n339) );
  OAI21_X1 U96 ( .B1(n444), .B2(n165), .A(n166), .ZN(n283) );
  OAI21_X1 U97 ( .B1(n444), .B2(n203), .A(n204), .ZN(n315) );
  OAI21_X1 U98 ( .B1(n444), .B2(n175), .A(n176), .ZN(n291) );
  OAI21_X1 U99 ( .B1(n444), .B2(n63), .A(n64), .ZN(n355) );
  NOR2_X1 U100 ( .A1(clr_delay), .A2(delay_timer[0]), .ZN(N108) );
  NOR2_X1 U101 ( .A1(addr_a[0]), .A2(clr_addr_a), .ZN(N89) );
  INV_X1 U102 ( .A(n399), .ZN(n400) );
  INV_X1 U103 ( .A(n395), .ZN(n396) );
  INV_X1 U104 ( .A(n216), .ZN(n217) );
  AND2_X1 U105 ( .A1(addr_a[0]), .A2(n12), .ZN(n52) );
  NAND2_X1 U106 ( .A1(addr_a[0]), .A2(addr_a[1]), .ZN(n225) );
  OAI21_X1 U107 ( .B1(n444), .B2(n128), .A(n129), .ZN(n251) );
  NAND2_X1 U108 ( .A1(n124), .A2(n128), .ZN(n129) );
  OAI21_X1 U109 ( .B1(n444), .B2(n110), .A(n111), .ZN(n235) );
  NAND2_X1 U110 ( .A1(n116), .A2(n110), .ZN(n111) );
  INV_X1 U111 ( .A(clr_addr_a), .ZN(n441) );
  OAI21_X1 U112 ( .B1(n444), .B2(n146), .A(n147), .ZN(n267) );
  NAND2_X1 U113 ( .A1(\a[14][7] ), .A2(n146), .ZN(n147) );
  OAI21_X1 U114 ( .B1(n444), .B2(n73), .A(n74), .ZN(n363) );
  OAI21_X1 U115 ( .B1(n444), .B2(n156), .A(n157), .ZN(n275) );
  OAI21_X1 U116 ( .B1(n444), .B2(n194), .A(n195), .ZN(n307) );
  OAI21_X1 U117 ( .B1(n444), .B2(n185), .A(n186), .ZN(n299) );
  OAI21_X1 U118 ( .B1(n444), .B2(n91), .A(n92), .ZN(n379) );
  OAI21_X1 U119 ( .B1(n444), .B2(n82), .A(n83), .ZN(n371) );
  OAI21_X1 U120 ( .B1(n32), .B2(n444), .A(n33), .ZN(n331) );
  AND2_X1 U121 ( .A1(n100), .A2(n10), .ZN(n72) );
  AND2_X1 U122 ( .A1(n174), .A2(n10), .ZN(n184) );
  AND2_X1 U123 ( .A1(N24), .A2(N25), .ZN(N116) );
  AND2_X1 U124 ( .A1(addr_a[2]), .A2(n100), .ZN(n42) );
  NOR2_X1 U125 ( .A1(clr_delay), .A2(n233), .ZN(N109) );
  XNOR2_X1 U126 ( .A(delay_timer[0]), .B(delay_timer[1]), .ZN(n233) );
  NOR2_X1 U127 ( .A1(clr_addr_y), .A2(n234), .ZN(N102) );
  XNOR2_X1 U128 ( .A(N25), .B(N24), .ZN(n234) );
  INV_X1 U129 ( .A(clr_delay), .ZN(n443) );
  NOR2_X1 U130 ( .A1(clr_addr_y), .A2(N24), .ZN(N101) );
  NOR2_X1 U131 ( .A1(clr_addr_x), .A2(n221), .ZN(N97) );
  XNOR2_X1 U132 ( .A(addr_x[1]), .B(addr_x[0]), .ZN(n221) );
  NOR2_X1 U133 ( .A1(clr_addr_x), .A2(addr_x[0]), .ZN(N96) );
  AND2_X1 U134 ( .A1(n174), .A2(addr_a[2]), .ZN(n155) );
  AND2_X1 U135 ( .A1(en_a), .A2(n9), .ZN(n100) );
  AND2_X1 U136 ( .A1(addr_a[3]), .A2(en_a), .ZN(n174) );
  INV_X1 U137 ( .A(n101), .ZN(n431) );
  MUX2_X1 U138 ( .A(\y[2][0] ), .B(\y[3][0] ), .S(n211), .Z(n168) );
  MUX2_X1 U139 ( .A(\y[0][0] ), .B(\y[1][0] ), .S(n211), .Z(n169) );
  MUX2_X1 U140 ( .A(n169), .B(n168), .S(N25), .Z(N83) );
  MUX2_X1 U141 ( .A(\y[2][1] ), .B(\y[3][1] ), .S(n211), .Z(n170) );
  MUX2_X1 U142 ( .A(\y[0][1] ), .B(\y[1][1] ), .S(n211), .Z(n171) );
  MUX2_X1 U143 ( .A(n171), .B(n170), .S(N25), .Z(N82) );
  MUX2_X1 U144 ( .A(\y[2][2] ), .B(\y[3][2] ), .S(n211), .Z(n172) );
  MUX2_X1 U145 ( .A(\y[0][2] ), .B(\y[1][2] ), .S(n211), .Z(n173) );
  MUX2_X1 U146 ( .A(n173), .B(n172), .S(N25), .Z(N81) );
  MUX2_X1 U147 ( .A(\y[2][3] ), .B(\y[3][3] ), .S(n211), .Z(n177) );
  MUX2_X1 U148 ( .A(\y[0][3] ), .B(\y[1][3] ), .S(n211), .Z(n178) );
  MUX2_X1 U149 ( .A(n178), .B(n177), .S(N25), .Z(N80) );
  MUX2_X1 U150 ( .A(\y[2][4] ), .B(\y[3][4] ), .S(n211), .Z(n179) );
  MUX2_X1 U151 ( .A(\y[0][4] ), .B(\y[1][4] ), .S(n211), .Z(n180) );
  MUX2_X1 U152 ( .A(n180), .B(n179), .S(N25), .Z(N79) );
  MUX2_X1 U153 ( .A(\y[2][5] ), .B(\y[3][5] ), .S(n211), .Z(n181) );
  MUX2_X1 U154 ( .A(\y[0][5] ), .B(\y[1][5] ), .S(n211), .Z(n182) );
  MUX2_X1 U155 ( .A(n182), .B(n181), .S(N25), .Z(N78) );
  MUX2_X1 U156 ( .A(\y[2][6] ), .B(\y[3][6] ), .S(N24), .Z(n183) );
  MUX2_X1 U157 ( .A(\y[0][6] ), .B(\y[1][6] ), .S(N24), .Z(n187) );
  MUX2_X1 U158 ( .A(n187), .B(n183), .S(N25), .Z(N77) );
  MUX2_X1 U159 ( .A(\y[2][7] ), .B(\y[3][7] ), .S(N24), .Z(n188) );
  MUX2_X1 U160 ( .A(\y[0][7] ), .B(\y[1][7] ), .S(n211), .Z(n189) );
  MUX2_X1 U161 ( .A(n189), .B(n188), .S(N25), .Z(N76) );
  MUX2_X1 U162 ( .A(\y[2][8] ), .B(\y[3][8] ), .S(n211), .Z(n190) );
  MUX2_X1 U163 ( .A(\y[0][8] ), .B(\y[1][8] ), .S(N24), .Z(n191) );
  MUX2_X1 U164 ( .A(n191), .B(n190), .S(N25), .Z(N75) );
  MUX2_X1 U165 ( .A(\y[2][9] ), .B(\y[3][9] ), .S(N24), .Z(n192) );
  MUX2_X1 U166 ( .A(\y[0][9] ), .B(\y[1][9] ), .S(N24), .Z(n193) );
  MUX2_X1 U167 ( .A(n193), .B(n192), .S(N25), .Z(N74) );
  MUX2_X1 U168 ( .A(\y[2][10] ), .B(\y[3][10] ), .S(N24), .Z(n196) );
  MUX2_X1 U169 ( .A(\y[0][10] ), .B(\y[1][10] ), .S(n211), .Z(n197) );
  MUX2_X1 U170 ( .A(n197), .B(n196), .S(N25), .Z(N73) );
  NAND2_X1 U171 ( .A1(n198), .A2(n199), .ZN(N72) );
  AOI22_X1 U172 ( .A1(\y[1][11] ), .A2(n1), .B1(\y[3][11] ), .B2(N116), .ZN(
        n199) );
  AOI22_X1 U173 ( .A1(\y[0][11] ), .A2(n2), .B1(\y[2][11] ), .B2(n3), .ZN(n198) );
  NAND2_X1 U174 ( .A1(n200), .A2(n201), .ZN(N71) );
  AOI22_X1 U175 ( .A1(\y[1][12] ), .A2(n1), .B1(\y[3][12] ), .B2(N116), .ZN(
        n201) );
  AOI22_X1 U176 ( .A1(\y[0][12] ), .A2(n2), .B1(\y[2][12] ), .B2(n3), .ZN(n200) );
  NAND2_X1 U177 ( .A1(n202), .A2(n205), .ZN(N70) );
  AOI22_X1 U178 ( .A1(\y[1][13] ), .A2(n1), .B1(\y[3][13] ), .B2(N116), .ZN(
        n205) );
  AOI22_X1 U179 ( .A1(\y[0][13] ), .A2(n2), .B1(\y[2][13] ), .B2(n3), .ZN(n202) );
  NAND2_X1 U180 ( .A1(n206), .A2(n207), .ZN(N69) );
  AOI22_X1 U181 ( .A1(\y[1][14] ), .A2(n1), .B1(\y[3][14] ), .B2(N116), .ZN(
        n207) );
  AOI22_X1 U182 ( .A1(\y[0][14] ), .A2(n2), .B1(\y[2][14] ), .B2(n3), .ZN(n206) );
  NAND2_X1 U183 ( .A1(n208), .A2(n209), .ZN(N68) );
  AOI22_X1 U184 ( .A1(\y[1][15] ), .A2(n1), .B1(\y[3][15] ), .B2(N116), .ZN(
        n209) );
  AOI22_X1 U185 ( .A1(\y[0][15] ), .A2(n2), .B1(\y[2][15] ), .B2(n3), .ZN(n208) );
  NAND2_X1 U186 ( .A1(\a[6][7] ), .A2(n32), .ZN(n33) );
  NAND2_X1 U187 ( .A1(\a[5][7] ), .A2(n43), .ZN(n44) );
  OAI21_X1 U188 ( .B1(n444), .B2(n53), .A(n54), .ZN(n347) );
  BUF_X4 U189 ( .A(\x[2][4] ), .Z(n214) );
  NAND2_X1 U190 ( .A1(\a[3][7] ), .A2(n63), .ZN(n64) );
  NAND2_X1 U191 ( .A1(\a[12][7] ), .A2(n165), .ZN(n166) );
  NAND2_X1 U192 ( .A1(\a[7][7] ), .A2(n212), .ZN(n213) );
  NAND2_X1 U193 ( .A1(\a[11][7] ), .A2(n175), .ZN(n176) );
  NAND2_X1 U194 ( .A1(\a[15][7] ), .A2(n137), .ZN(n138) );
  INV_X2 U195 ( .A(n387), .ZN(n388) );
  INV_X2 U196 ( .A(n389), .ZN(n390) );
  NAND2_X1 U197 ( .A1(\a[10][7] ), .A2(n185), .ZN(n186) );
  NAND2_X1 U198 ( .A1(\a[0][7] ), .A2(n91), .ZN(n92) );
  NAND2_X1 U199 ( .A1(\a[1][7] ), .A2(n82), .ZN(n83) );
  NAND2_X1 U200 ( .A1(\a[13][7] ), .A2(n156), .ZN(n157) );
  INV_X2 U201 ( .A(n393), .ZN(n394) );
  NAND2_X1 U202 ( .A1(\a[2][7] ), .A2(n73), .ZN(n74) );
  NAND2_X1 U203 ( .A1(\a[8][7] ), .A2(n203), .ZN(n204) );
  NAND2_X1 U204 ( .A1(n132), .A2(n194), .ZN(n195) );
  INV_X2 U205 ( .A(n401), .ZN(n402) );
  NAND2_X1 U206 ( .A1(\a[4][7] ), .A2(n53), .ZN(n54) );
  INV_X2 U207 ( .A(n403), .ZN(n404) );
  INV_X2 U208 ( .A(n407), .ZN(n408) );
  INV_X1 U209 ( .A(n409), .ZN(n410) );
  NAND2_X1 U210 ( .A1(n122), .A2(n119), .ZN(n120) );
  AOI22_X1 U211 ( .A1(data_in[7]), .A2(n439), .B1(n102), .B2(n81), .ZN(n101)
         );
  NAND2_X1 U212 ( .A1(en_a), .A2(N114), .ZN(n137) );
  INV_X1 U213 ( .A(n137), .ZN(n411) );
  MUX2_X1 U214 ( .A(\a[15][6] ), .B(data_in[6]), .S(n411), .Z(n260) );
  MUX2_X1 U215 ( .A(\a[15][5] ), .B(data_in[5]), .S(n411), .Z(n261) );
  MUX2_X1 U216 ( .A(\a[15][4] ), .B(data_in[4]), .S(n411), .Z(n262) );
  MUX2_X1 U217 ( .A(n150), .B(data_in[3]), .S(n411), .Z(n263) );
  MUX2_X1 U218 ( .A(\a[15][2] ), .B(data_in[2]), .S(n411), .Z(n264) );
  MUX2_X1 U219 ( .A(\a[15][1] ), .B(data_in[1]), .S(n411), .Z(n265) );
  MUX2_X1 U220 ( .A(\a[15][0] ), .B(data_in[0]), .S(n411), .Z(n266) );
  NAND2_X1 U221 ( .A1(n155), .A2(n41), .ZN(n146) );
  INV_X1 U222 ( .A(n146), .ZN(n412) );
  MUX2_X1 U223 ( .A(\a[14][6] ), .B(data_in[6]), .S(n412), .Z(n268) );
  MUX2_X1 U224 ( .A(\a[14][5] ), .B(data_in[5]), .S(n412), .Z(n269) );
  MUX2_X1 U225 ( .A(\a[14][4] ), .B(data_in[4]), .S(n412), .Z(n270) );
  MUX2_X1 U226 ( .A(\a[14][3] ), .B(data_in[3]), .S(n412), .Z(n271) );
  MUX2_X1 U227 ( .A(n13), .B(data_in[2]), .S(n412), .Z(n272) );
  MUX2_X1 U228 ( .A(n219), .B(data_in[1]), .S(n412), .Z(n273) );
  MUX2_X1 U229 ( .A(\a[14][0] ), .B(data_in[0]), .S(n412), .Z(n274) );
  NAND2_X1 U230 ( .A1(n155), .A2(n52), .ZN(n156) );
  INV_X1 U231 ( .A(n156), .ZN(n413) );
  MUX2_X1 U232 ( .A(\a[13][6] ), .B(data_in[6]), .S(n413), .Z(n276) );
  MUX2_X1 U233 ( .A(\a[13][5] ), .B(data_in[5]), .S(n413), .Z(n277) );
  MUX2_X1 U234 ( .A(\a[13][4] ), .B(data_in[4]), .S(n413), .Z(n278) );
  MUX2_X1 U235 ( .A(\a[13][3] ), .B(data_in[3]), .S(n413), .Z(n279) );
  MUX2_X1 U236 ( .A(\a[13][2] ), .B(data_in[2]), .S(n413), .Z(n280) );
  MUX2_X1 U237 ( .A(\a[13][1] ), .B(data_in[1]), .S(n413), .Z(n281) );
  MUX2_X1 U238 ( .A(\a[13][0] ), .B(data_in[0]), .S(n413), .Z(n282) );
  NAND2_X1 U239 ( .A1(n155), .A2(n62), .ZN(n165) );
  INV_X1 U240 ( .A(n165), .ZN(n414) );
  MUX2_X1 U241 ( .A(\a[12][6] ), .B(data_in[6]), .S(n414), .Z(n284) );
  MUX2_X1 U242 ( .A(\a[12][5] ), .B(data_in[5]), .S(n414), .Z(n285) );
  MUX2_X1 U243 ( .A(\a[12][4] ), .B(data_in[4]), .S(n414), .Z(n286) );
  MUX2_X1 U244 ( .A(n8), .B(data_in[3]), .S(n414), .Z(n287) );
  MUX2_X1 U245 ( .A(\a[12][2] ), .B(data_in[2]), .S(n414), .Z(n288) );
  MUX2_X1 U246 ( .A(\a[12][1] ), .B(data_in[1]), .S(n414), .Z(n289) );
  MUX2_X1 U247 ( .A(\a[12][0] ), .B(data_in[0]), .S(n414), .Z(n290) );
  NAND2_X1 U248 ( .A1(en_x), .A2(N115), .ZN(n102) );
  INV_X1 U249 ( .A(n102), .ZN(n439) );
  MUX2_X1 U250 ( .A(n70), .B(data_in[6]), .S(n439), .Z(n432) );
  MUX2_X1 U251 ( .A(\x[3][5] ), .B(data_in[5]), .S(n439), .Z(n433) );
  MUX2_X1 U252 ( .A(\x[3][4] ), .B(data_in[4]), .S(n439), .Z(n434) );
  MUX2_X1 U253 ( .A(n55), .B(data_in[3]), .S(n439), .Z(n435) );
  MUX2_X1 U254 ( .A(n97), .B(data_in[2]), .S(n439), .Z(n436) );
  MUX2_X1 U255 ( .A(n217), .B(data_in[1]), .S(n439), .Z(n437) );
  MUX2_X1 U256 ( .A(\x[3][0] ), .B(data_in[0]), .S(n439), .Z(n438) );
  NAND3_X1 U257 ( .A1(addr_x[1]), .A2(n16), .A3(en_x), .ZN(n110) );
  INV_X1 U258 ( .A(n110), .ZN(n415) );
  MUX2_X1 U259 ( .A(n40), .B(data_in[6]), .S(n415), .Z(n236) );
  MUX2_X1 U260 ( .A(n48), .B(data_in[5]), .S(n415), .Z(n237) );
  MUX2_X1 U261 ( .A(n214), .B(data_in[4]), .S(n415), .Z(n238) );
  MUX2_X1 U262 ( .A(n89), .B(data_in[3]), .S(n415), .Z(n239) );
  MUX2_X1 U263 ( .A(n215), .B(data_in[2]), .S(n415), .Z(n240) );
  MUX2_X1 U264 ( .A(n159), .B(data_in[1]), .S(n415), .Z(n241) );
  MUX2_X1 U265 ( .A(n36), .B(data_in[0]), .S(n415), .Z(n242) );
  NAND3_X1 U266 ( .A1(addr_x[0]), .A2(n15), .A3(en_x), .ZN(n119) );
  INV_X1 U267 ( .A(n119), .ZN(n416) );
  MUX2_X1 U268 ( .A(n75), .B(data_in[6]), .S(n416), .Z(n244) );
  MUX2_X1 U269 ( .A(n59), .B(data_in[5]), .S(n416), .Z(n245) );
  MUX2_X1 U270 ( .A(n38), .B(data_in[4]), .S(n416), .Z(n246) );
  MUX2_X1 U271 ( .A(n396), .B(data_in[3]), .S(n416), .Z(n247) );
  MUX2_X1 U272 ( .A(n66), .B(data_in[2]), .S(n416), .Z(n248) );
  MUX2_X1 U273 ( .A(n130), .B(data_in[1]), .S(n416), .Z(n249) );
  MUX2_X1 U274 ( .A(n24), .B(data_in[0]), .S(n416), .Z(n250) );
  NAND3_X1 U275 ( .A1(n15), .A2(n16), .A3(en_x), .ZN(n128) );
  INV_X1 U276 ( .A(n128), .ZN(n417) );
  MUX2_X1 U277 ( .A(n85), .B(data_in[6]), .S(n417), .Z(n252) );
  MUX2_X1 U278 ( .A(n61), .B(data_in[5]), .S(n417), .Z(n253) );
  MUX2_X1 U279 ( .A(n126), .B(data_in[4]), .S(n417), .Z(n254) );
  MUX2_X1 U280 ( .A(\x[0][3] ), .B(data_in[3]), .S(n417), .Z(n255) );
  MUX2_X1 U281 ( .A(n87), .B(data_in[2]), .S(n417), .Z(n256) );
  MUX2_X1 U282 ( .A(n400), .B(data_in[1]), .S(n417), .Z(n257) );
  MUX2_X1 U283 ( .A(\x[0][0] ), .B(data_in[0]), .S(n417), .Z(n258) );
  INV_X1 U284 ( .A(n225), .ZN(n430) );
  NAND2_X1 U285 ( .A1(n184), .A2(n430), .ZN(n175) );
  INV_X1 U286 ( .A(n175), .ZN(n418) );
  MUX2_X1 U287 ( .A(\a[11][6] ), .B(data_in[6]), .S(n418), .Z(n292) );
  MUX2_X1 U288 ( .A(\a[11][5] ), .B(data_in[5]), .S(n418), .Z(n293) );
  MUX2_X1 U289 ( .A(\a[11][4] ), .B(data_in[4]), .S(n418), .Z(n294) );
  MUX2_X1 U290 ( .A(n106), .B(data_in[3]), .S(n418), .Z(n295) );
  MUX2_X1 U291 ( .A(\a[11][2] ), .B(data_in[2]), .S(n418), .Z(n296) );
  MUX2_X1 U292 ( .A(n112), .B(data_in[1]), .S(n418), .Z(n297) );
  MUX2_X1 U293 ( .A(\a[11][0] ), .B(data_in[0]), .S(n418), .Z(n298) );
  NAND2_X1 U294 ( .A1(n184), .A2(n41), .ZN(n185) );
  INV_X1 U295 ( .A(n185), .ZN(n419) );
  MUX2_X1 U296 ( .A(\a[10][6] ), .B(data_in[6]), .S(n419), .Z(n300) );
  MUX2_X1 U297 ( .A(\a[10][5] ), .B(data_in[5]), .S(n419), .Z(n301) );
  MUX2_X1 U298 ( .A(\a[10][4] ), .B(data_in[4]), .S(n419), .Z(n302) );
  MUX2_X1 U299 ( .A(\a[10][3] ), .B(data_in[3]), .S(n419), .Z(n303) );
  MUX2_X1 U300 ( .A(\a[10][2] ), .B(data_in[2]), .S(n419), .Z(n304) );
  MUX2_X1 U301 ( .A(n34), .B(data_in[1]), .S(n419), .Z(n305) );
  MUX2_X1 U302 ( .A(\a[10][0] ), .B(data_in[0]), .S(n419), .Z(n306) );
  NAND2_X1 U303 ( .A1(n184), .A2(n52), .ZN(n194) );
  INV_X1 U304 ( .A(n194), .ZN(n420) );
  MUX2_X1 U305 ( .A(n79), .B(data_in[6]), .S(n420), .Z(n308) );
  MUX2_X1 U306 ( .A(\a[9][5] ), .B(data_in[5]), .S(n420), .Z(n309) );
  MUX2_X1 U307 ( .A(\a[9][4] ), .B(data_in[4]), .S(n420), .Z(n310) );
  MUX2_X1 U308 ( .A(n392), .B(data_in[3]), .S(n420), .Z(n311) );
  MUX2_X1 U309 ( .A(\a[9][2] ), .B(data_in[2]), .S(n420), .Z(n312) );
  MUX2_X1 U310 ( .A(n93), .B(data_in[1]), .S(n420), .Z(n313) );
  MUX2_X1 U311 ( .A(\a[9][0] ), .B(data_in[0]), .S(n420), .Z(n314) );
  NAND2_X1 U312 ( .A1(n184), .A2(n62), .ZN(n203) );
  INV_X1 U313 ( .A(n203), .ZN(n421) );
  MUX2_X1 U314 ( .A(n28), .B(data_in[6]), .S(n421), .Z(n316) );
  MUX2_X1 U315 ( .A(\a[8][5] ), .B(data_in[5]), .S(n421), .Z(n317) );
  MUX2_X1 U316 ( .A(\a[8][4] ), .B(data_in[4]), .S(n421), .Z(n318) );
  MUX2_X1 U317 ( .A(n30), .B(data_in[3]), .S(n421), .Z(n319) );
  MUX2_X1 U318 ( .A(n50), .B(data_in[2]), .S(n421), .Z(n320) );
  MUX2_X1 U319 ( .A(n104), .B(data_in[1]), .S(n421), .Z(n321) );
  MUX2_X1 U320 ( .A(\a[8][0] ), .B(data_in[0]), .S(n421), .Z(n322) );
  NAND2_X1 U321 ( .A1(n42), .A2(n430), .ZN(n212) );
  INV_X1 U322 ( .A(n212), .ZN(n422) );
  MUX2_X1 U323 ( .A(\a[7][6] ), .B(data_in[6]), .S(n422), .Z(n324) );
  MUX2_X1 U324 ( .A(n161), .B(data_in[5]), .S(n422), .Z(n325) );
  MUX2_X1 U325 ( .A(\a[7][4] ), .B(data_in[4]), .S(n422), .Z(n326) );
  MUX2_X1 U326 ( .A(\a[7][3] ), .B(data_in[3]), .S(n422), .Z(n327) );
  MUX2_X1 U327 ( .A(\a[7][2] ), .B(data_in[2]), .S(n422), .Z(n328) );
  MUX2_X1 U328 ( .A(\a[7][1] ), .B(data_in[1]), .S(n422), .Z(n329) );
  MUX2_X1 U329 ( .A(\a[7][0] ), .B(data_in[0]), .S(n422), .Z(n330) );
  NAND2_X1 U330 ( .A1(n42), .A2(n41), .ZN(n32) );
  INV_X1 U331 ( .A(n32), .ZN(n423) );
  MUX2_X1 U332 ( .A(\a[6][6] ), .B(data_in[6]), .S(n423), .Z(n332) );
  MUX2_X1 U333 ( .A(\a[6][5] ), .B(data_in[5]), .S(n423), .Z(n333) );
  MUX2_X1 U334 ( .A(\a[6][4] ), .B(data_in[4]), .S(n423), .Z(n334) );
  MUX2_X1 U335 ( .A(\a[6][3] ), .B(data_in[3]), .S(n423), .Z(n335) );
  MUX2_X1 U336 ( .A(\a[6][2] ), .B(data_in[2]), .S(n423), .Z(n336) );
  MUX2_X1 U337 ( .A(\a[6][1] ), .B(data_in[1]), .S(n423), .Z(n337) );
  MUX2_X1 U338 ( .A(\a[6][0] ), .B(data_in[0]), .S(n423), .Z(n338) );
  NAND2_X1 U339 ( .A1(n42), .A2(n52), .ZN(n43) );
  INV_X1 U340 ( .A(n43), .ZN(n424) );
  MUX2_X1 U341 ( .A(\a[5][6] ), .B(data_in[6]), .S(n424), .Z(n340) );
  MUX2_X1 U342 ( .A(\a[5][5] ), .B(data_in[5]), .S(n424), .Z(n341) );
  MUX2_X1 U343 ( .A(\a[5][4] ), .B(data_in[4]), .S(n424), .Z(n342) );
  MUX2_X1 U344 ( .A(n134), .B(data_in[3]), .S(n424), .Z(n343) );
  MUX2_X1 U345 ( .A(\a[5][2] ), .B(data_in[2]), .S(n424), .Z(n344) );
  MUX2_X1 U346 ( .A(\a[5][1] ), .B(data_in[1]), .S(n424), .Z(n345) );
  MUX2_X1 U347 ( .A(\a[5][0] ), .B(data_in[0]), .S(n424), .Z(n346) );
  NAND2_X1 U348 ( .A1(n42), .A2(n62), .ZN(n53) );
  INV_X1 U349 ( .A(n53), .ZN(n425) );
  MUX2_X1 U350 ( .A(\a[4][6] ), .B(data_in[6]), .S(n425), .Z(n348) );
  MUX2_X1 U351 ( .A(n144), .B(data_in[5]), .S(n425), .Z(n349) );
  MUX2_X1 U352 ( .A(\a[4][4] ), .B(data_in[4]), .S(n425), .Z(n350) );
  MUX2_X1 U353 ( .A(\a[4][3] ), .B(data_in[3]), .S(n425), .Z(n351) );
  MUX2_X1 U354 ( .A(n22), .B(data_in[2]), .S(n425), .Z(n352) );
  MUX2_X1 U355 ( .A(n398), .B(data_in[1]), .S(n425), .Z(n353) );
  MUX2_X1 U356 ( .A(\a[4][0] ), .B(data_in[0]), .S(n425), .Z(n354) );
  NAND2_X1 U357 ( .A1(n72), .A2(n430), .ZN(n63) );
  INV_X1 U358 ( .A(n63), .ZN(n426) );
  MUX2_X1 U359 ( .A(\a[3][6] ), .B(data_in[6]), .S(n426), .Z(n356) );
  MUX2_X1 U360 ( .A(\a[3][5] ), .B(data_in[5]), .S(n426), .Z(n357) );
  MUX2_X1 U361 ( .A(\a[3][4] ), .B(data_in[4]), .S(n426), .Z(n358) );
  MUX2_X1 U362 ( .A(\a[3][3] ), .B(data_in[3]), .S(n426), .Z(n359) );
  MUX2_X1 U363 ( .A(\a[3][2] ), .B(data_in[2]), .S(n426), .Z(n360) );
  MUX2_X1 U364 ( .A(n77), .B(data_in[1]), .S(n426), .Z(n361) );
  MUX2_X1 U365 ( .A(\a[3][0] ), .B(data_in[0]), .S(n426), .Z(n362) );
  NAND2_X1 U366 ( .A1(n41), .A2(n72), .ZN(n73) );
  INV_X1 U367 ( .A(n73), .ZN(n427) );
  MUX2_X1 U368 ( .A(\a[2][6] ), .B(data_in[6]), .S(n427), .Z(n364) );
  MUX2_X1 U369 ( .A(\a[2][5] ), .B(data_in[5]), .S(n427), .Z(n365) );
  MUX2_X1 U370 ( .A(\a[2][4] ), .B(data_in[4]), .S(n427), .Z(n366) );
  MUX2_X1 U371 ( .A(\a[2][3] ), .B(data_in[3]), .S(n427), .Z(n367) );
  MUX2_X1 U372 ( .A(\a[2][2] ), .B(data_in[2]), .S(n427), .Z(n368) );
  MUX2_X1 U373 ( .A(\a[2][1] ), .B(data_in[1]), .S(n427), .Z(n369) );
  MUX2_X1 U374 ( .A(\a[2][0] ), .B(data_in[0]), .S(n427), .Z(n370) );
  NAND2_X1 U375 ( .A1(n52), .A2(n72), .ZN(n82) );
  INV_X1 U376 ( .A(n82), .ZN(n428) );
  MUX2_X1 U377 ( .A(n118), .B(data_in[6]), .S(n428), .Z(n372) );
  MUX2_X1 U378 ( .A(n57), .B(data_in[5]), .S(n428), .Z(n373) );
  MUX2_X1 U379 ( .A(\a[1][4] ), .B(data_in[4]), .S(n428), .Z(n374) );
  MUX2_X1 U380 ( .A(n99), .B(data_in[3]), .S(n428), .Z(n375) );
  MUX2_X1 U381 ( .A(\a[1][2] ), .B(data_in[2]), .S(n428), .Z(n376) );
  MUX2_X1 U382 ( .A(n410), .B(data_in[1]), .S(n428), .Z(n377) );
  MUX2_X1 U383 ( .A(\a[1][0] ), .B(data_in[0]), .S(n428), .Z(n378) );
  NAND2_X1 U384 ( .A1(n72), .A2(n62), .ZN(n91) );
  INV_X1 U385 ( .A(n91), .ZN(n429) );
  MUX2_X1 U386 ( .A(\a[0][6] ), .B(data_in[6]), .S(n429), .Z(n380) );
  MUX2_X1 U387 ( .A(\a[0][5] ), .B(data_in[5]), .S(n429), .Z(n381) );
  MUX2_X1 U388 ( .A(n17), .B(data_in[4]), .S(n429), .Z(n382) );
  MUX2_X1 U389 ( .A(n6), .B(data_in[3]), .S(n429), .Z(n383) );
  MUX2_X1 U390 ( .A(\a[0][2] ), .B(data_in[2]), .S(n429), .Z(n384) );
  MUX2_X1 U391 ( .A(\a[0][1] ), .B(data_in[1]), .S(n429), .Z(n385) );
  MUX2_X1 U392 ( .A(\a[0][0] ), .B(data_in[0]), .S(n429), .Z(n386) );
endmodule


module control_DELAY2 ( clk, reset, start, done, en_a, en_x, en_y, clr_addr_a, 
        clr_addr_x, clr_addr_y, clr_delay, of_a, of_x, of_y, of_delay );
  input clk, reset, start, of_a, of_x, of_y, of_delay;
  output done, en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay;
  wire   \in_state[1] , n1, n7, n8, n12, n14, n15, n16, n17, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n2, n3, n4, n5, n6, n9,
         n10, n11, n13, n18, n19, n20, n21;
  wire   [1:0] out_state;
  assign en_y = 1'b0;

  DFF_X1 \in_state_reg[0]  ( .D(n61), .CK(clk), .QN(n8) );
  DFF_X1 \in_state_reg[1]  ( .D(n60), .CK(clk), .Q(\in_state[1] ), .QN(n7) );
  DFF_X1 \out_state_reg[0]  ( .D(n59), .CK(clk), .Q(out_state[0]), .QN(n14) );
  DFF_X1 \out_state_reg[1]  ( .D(n58), .CK(clk), .Q(out_state[1]), .QN(n12) );
  DFF_X1 done_reg ( .D(n57), .CK(clk), .Q(done), .QN(n1) );
  DFF_X1 en_a_reg ( .D(n56), .CK(clk), .Q(en_a) );
  DFF_X1 en_x_reg ( .D(n55), .CK(clk), .Q(en_x) );
  DFF_X1 clr_addr_a_reg ( .D(n54), .CK(clk), .Q(clr_addr_a), .QN(n15) );
  DFF_X1 clr_addr_x_reg ( .D(n53), .CK(clk), .Q(clr_addr_x), .QN(n16) );
  DFF_X1 clr_addr_y_reg ( .D(n52), .CK(clk), .Q(clr_addr_y), .QN(n17) );
  DFF_X1 clr_delay_reg ( .D(n6), .CK(clk), .Q(clr_delay) );
  NAND3_X1 U51 ( .A1(of_delay), .A2(n12), .A3(out_state[0]), .ZN(n28) );
  NAND3_X1 U52 ( .A1(n29), .A2(n20), .A3(n33), .ZN(n35) );
  NAND3_X1 U53 ( .A1(n12), .A2(n20), .A3(out_state[0]), .ZN(n43) );
  NAND3_X1 U54 ( .A1(n8), .A2(n14), .A3(n45), .ZN(n46) );
  NAND3_X1 U55 ( .A1(n48), .A2(n20), .A3(n33), .ZN(n49) );
  NAND3_X1 U56 ( .A1(n48), .A2(n20), .A3(n51), .ZN(n50) );
  INV_X1 U4 ( .A(n29), .ZN(n5) );
  INV_X1 U5 ( .A(n31), .ZN(n2) );
  OAI21_X1 U6 ( .B1(n21), .B2(n40), .A(n5), .ZN(n48) );
  OAI21_X1 U7 ( .B1(n38), .B2(n21), .A(n39), .ZN(n31) );
  AOI21_X1 U8 ( .B1(n4), .B2(of_x), .A(n3), .ZN(n38) );
  OAI21_X1 U9 ( .B1(n18), .B2(n41), .A(n39), .ZN(n29) );
  INV_X1 U10 ( .A(n41), .ZN(n4) );
  INV_X1 U11 ( .A(of_delay), .ZN(n19) );
  INV_X1 U12 ( .A(n40), .ZN(n3) );
  INV_X1 U13 ( .A(of_x), .ZN(n18) );
  NOR2_X1 U14 ( .A1(n8), .A2(\in_state[1] ), .ZN(n33) );
  AOI21_X1 U15 ( .B1(out_state[0]), .B2(out_state[1]), .A(reset), .ZN(n26) );
  AOI21_X1 U16 ( .B1(n33), .B2(of_a), .A(reset), .ZN(n39) );
  OAI22_X1 U17 ( .A1(n42), .A2(n1), .B1(n10), .B2(n43), .ZN(n57) );
  INV_X1 U18 ( .A(n42), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n19), .B2(n14), .A(n26), .ZN(n42) );
  OAI22_X1 U20 ( .A1(n25), .A2(n17), .B1(n11), .B2(n26), .ZN(n52) );
  INV_X1 U21 ( .A(n25), .ZN(n11) );
  OAI21_X1 U22 ( .B1(n27), .B2(n12), .A(n13), .ZN(n25) );
  INV_X1 U23 ( .A(n24), .ZN(n13) );
  OAI22_X1 U24 ( .A1(n29), .A2(n16), .B1(n5), .B2(n30), .ZN(n53) );
  NOR2_X1 U25 ( .A1(n4), .A2(reset), .ZN(n30) );
  OAI22_X1 U26 ( .A1(n31), .A2(n15), .B1(n2), .B2(n32), .ZN(n54) );
  NOR2_X1 U27 ( .A1(n33), .A2(reset), .ZN(n32) );
  NAND2_X1 U28 ( .A1(n8), .A2(n7), .ZN(n40) );
  NOR2_X1 U29 ( .A1(n18), .A2(n7), .ZN(n45) );
  NAND2_X1 U30 ( .A1(\in_state[1] ), .A2(n8), .ZN(n41) );
  AOI21_X1 U31 ( .B1(n9), .B2(n46), .A(reset), .ZN(n59) );
  INV_X1 U32 ( .A(n47), .ZN(n9) );
  AOI21_X1 U33 ( .B1(of_y), .B2(out_state[1]), .A(n14), .ZN(n47) );
  OAI21_X1 U34 ( .B1(n8), .B2(n48), .A(n50), .ZN(n61) );
  OAI21_X1 U35 ( .B1(n41), .B2(n21), .A(n40), .ZN(n51) );
  NAND2_X1 U36 ( .A1(n45), .A2(n8), .ZN(n23) );
  OAI21_X1 U37 ( .B1(n7), .B2(n48), .A(n49), .ZN(n60) );
  NAND2_X1 U38 ( .A1(n20), .A2(n28), .ZN(n24) );
  OAI21_X1 U39 ( .B1(n19), .B2(n43), .A(n44), .ZN(n58) );
  NAND4_X1 U40 ( .A1(out_state[1]), .A2(n27), .A3(n23), .A4(n20), .ZN(n44) );
  NAND2_X1 U41 ( .A1(of_y), .A2(out_state[0]), .ZN(n27) );
  NAND2_X1 U42 ( .A1(n34), .A2(n35), .ZN(n55) );
  NAND2_X1 U43 ( .A1(en_x), .A2(n5), .ZN(n34) );
  NAND2_X1 U44 ( .A1(n36), .A2(n37), .ZN(n56) );
  OAI211_X1 U45 ( .C1(n3), .C2(n4), .A(n31), .B(n20), .ZN(n37) );
  NAND2_X1 U46 ( .A1(en_a), .A2(n2), .ZN(n36) );
  INV_X1 U47 ( .A(n22), .ZN(n6) );
  AOI21_X1 U48 ( .B1(n23), .B2(clr_delay), .A(n24), .ZN(n22) );
  INV_X1 U49 ( .A(reset), .ZN(n20) );
  INV_X1 U50 ( .A(start), .ZN(n21) );
endmodule


module mvm4_part3 ( clk, reset, start, done, data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, start;
  output done;
  wire   en_a, en_x, clr_addr_a, clr_addr_x, clr_addr_y, clr_delay, of_a, of_x,
         of_y, of_delay;

  data_path_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_INTERREG1_DELAY2 datapath ( 
        .clk(clk), .en_a(en_a), .en_x(en_x), .en_y(1'b0), .clr_addr_a(
        clr_addr_a), .clr_addr_x(clr_addr_x), .clr_addr_y(clr_addr_y), 
        .clr_delay(clr_delay), .of_a(of_a), .of_x(of_x), .of_y(of_y), 
        .of_delay(of_delay), .data_in(data_in), .data_out(data_out) );
  control_DELAY2 ctrl ( .clk(clk), .reset(reset), .start(start), .done(done), 
        .en_a(en_a), .en_x(en_x), .clr_addr_a(clr_addr_a), .clr_addr_x(
        clr_addr_x), .clr_addr_y(clr_addr_y), .clr_delay(clr_delay), .of_a(
        of_a), .of_x(of_x), .of_y(of_y), .of_delay(of_delay) );
endmodule

