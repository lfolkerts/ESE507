
module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n12, n13, n14, n15, n16, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50,
         n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102, n103,
         n104, n105, n108, n109, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n153, n154, n155, n157, n158, n160, n161, n163, n164, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n245, n246, n247, n248, n250, n251, n252,
         n253, n254, n255, n256, n258, n259, n260, n261, n262, n263, n264,
         n265, n273, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n368, n369, n370, n371, n372, n373, n374;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n324), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  CLKBUF_X1 U268 ( .A(n263), .Z(n303) );
  CLKBUF_X2 U269 ( .A(n255), .Z(n372) );
  CLKBUF_X1 U270 ( .A(n73), .Z(n304) );
  BUF_X1 U271 ( .A(n222), .Z(n305) );
  CLKBUF_X1 U272 ( .A(n372), .Z(n306) );
  OR2_X1 U273 ( .A1(n344), .A2(n164), .ZN(n307) );
  OR2_X1 U274 ( .A1(n344), .A2(n164), .ZN(n308) );
  OR2_X1 U275 ( .A1(n344), .A2(n164), .ZN(n253) );
  NOR2_X1 U276 ( .A1(n64), .A2(n61), .ZN(n309) );
  NOR2_X2 U277 ( .A1(n121), .A2(n124), .ZN(n61) );
  OAI21_X2 U278 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  XNOR2_X1 U279 ( .A(n265), .B(a[2]), .ZN(n310) );
  AOI21_X1 U280 ( .B1(n366), .B2(n83), .A(n334), .ZN(n311) );
  OAI21_X1 U281 ( .B1(n78), .B2(n76), .A(n77), .ZN(n312) );
  BUF_X2 U282 ( .A(n368), .Z(n348) );
  XOR2_X1 U283 ( .A(n368), .B(a[2]), .Z(n313) );
  XOR2_X1 U284 ( .A(n368), .B(a[2]), .Z(n248) );
  NAND2_X1 U285 ( .A1(a[6]), .A2(n315), .ZN(n316) );
  NAND2_X1 U286 ( .A1(n314), .A2(n262), .ZN(n317) );
  NAND2_X1 U287 ( .A1(n316), .A2(n317), .ZN(n246) );
  INV_X1 U288 ( .A(a[6]), .ZN(n314) );
  INV_X1 U289 ( .A(n262), .ZN(n315) );
  CLKBUF_X1 U290 ( .A(n265), .Z(n318) );
  BUF_X2 U291 ( .A(n264), .Z(n368) );
  OR2_X1 U292 ( .A1(n147), .A2(n150), .ZN(n319) );
  INV_X1 U293 ( .A(n75), .ZN(n320) );
  CLKBUF_X1 U294 ( .A(n83), .Z(n321) );
  CLKBUF_X1 U295 ( .A(n263), .Z(n322) );
  BUF_X2 U296 ( .A(n245), .Z(n323) );
  OAI22_X1 U297 ( .A1(n339), .A2(n221), .B1(n220), .B2(n373), .ZN(n324) );
  OAI21_X1 U298 ( .B1(n61), .B2(n65), .A(n62), .ZN(n325) );
  INV_X1 U299 ( .A(n161), .ZN(n326) );
  BUF_X2 U300 ( .A(n350), .Z(n373) );
  XNOR2_X1 U301 ( .A(n133), .B(n327), .ZN(n131) );
  XNOR2_X1 U302 ( .A(n138), .B(n135), .ZN(n327) );
  CLKBUF_X1 U303 ( .A(n78), .Z(n328) );
  BUF_X2 U304 ( .A(n368), .Z(n347) );
  NAND2_X1 U305 ( .A1(n356), .A2(n357), .ZN(n329) );
  INV_X1 U306 ( .A(n261), .ZN(n330) );
  BUF_X1 U307 ( .A(n255), .Z(n371) );
  INV_X1 U308 ( .A(n64), .ZN(n103) );
  AND2_X1 U309 ( .A1(n335), .A2(n199), .ZN(n331) );
  OR2_X1 U310 ( .A1(n201), .A2(n169), .ZN(n332) );
  INV_X1 U311 ( .A(n355), .ZN(n333) );
  INV_X1 U312 ( .A(n72), .ZN(n105) );
  AND2_X1 U313 ( .A1(n147), .A2(n150), .ZN(n334) );
  XOR2_X1 U314 ( .A(n192), .B(n199), .Z(n153) );
  CLKBUF_X1 U315 ( .A(n192), .Z(n335) );
  NAND2_X1 U316 ( .A1(n133), .A2(n138), .ZN(n336) );
  NAND2_X1 U317 ( .A1(n133), .A2(n135), .ZN(n337) );
  NAND2_X1 U318 ( .A1(n138), .A2(n135), .ZN(n338) );
  NAND3_X1 U319 ( .A1(n336), .A2(n337), .A3(n338), .ZN(n130) );
  NAND2_X1 U320 ( .A1(n256), .A2(n313), .ZN(n339) );
  XOR2_X1 U321 ( .A(n148), .B(n183), .Z(n340) );
  XOR2_X1 U322 ( .A(n145), .B(n340), .Z(n143) );
  NAND2_X1 U323 ( .A1(n145), .A2(n148), .ZN(n341) );
  NAND2_X1 U324 ( .A1(n145), .A2(n183), .ZN(n342) );
  NAND2_X1 U325 ( .A1(n148), .A2(n183), .ZN(n343) );
  NAND3_X1 U326 ( .A1(n341), .A2(n342), .A3(n343), .ZN(n142) );
  XNOR2_X1 U327 ( .A(n265), .B(n164), .ZN(n344) );
  INV_X1 U328 ( .A(n164), .ZN(n273) );
  BUF_X1 U329 ( .A(n1), .Z(n369) );
  INV_X1 U330 ( .A(n259), .ZN(n345) );
  BUF_X2 U331 ( .A(n245), .Z(n374) );
  OR2_X1 U332 ( .A1(n143), .A2(n146), .ZN(n346) );
  NOR2_X1 U333 ( .A1(n131), .A2(n136), .ZN(n349) );
  NOR2_X1 U334 ( .A1(n131), .A2(n136), .ZN(n69) );
  XNOR2_X1 U335 ( .A(n265), .B(a[2]), .ZN(n350) );
  BUF_X2 U336 ( .A(n362), .Z(n351) );
  XNOR2_X1 U337 ( .A(n263), .B(a[6]), .ZN(n362) );
  NAND2_X1 U338 ( .A1(n329), .A2(n371), .ZN(n352) );
  NAND2_X1 U339 ( .A1(n329), .A2(n371), .ZN(n353) );
  NAND2_X1 U340 ( .A1(n247), .A2(n371), .ZN(n251) );
  NAND2_X1 U341 ( .A1(n263), .A2(n355), .ZN(n356) );
  NAND2_X1 U342 ( .A1(n354), .A2(n333), .ZN(n357) );
  NAND2_X1 U343 ( .A1(n356), .A2(n357), .ZN(n247) );
  INV_X1 U344 ( .A(n263), .ZN(n354) );
  INV_X1 U345 ( .A(a[4]), .ZN(n355) );
  NAND2_X1 U346 ( .A1(n313), .A2(n310), .ZN(n358) );
  NAND2_X1 U347 ( .A1(n248), .A2(n256), .ZN(n359) );
  NAND2_X1 U348 ( .A1(n246), .A2(n254), .ZN(n360) );
  NAND2_X1 U349 ( .A1(n246), .A2(n254), .ZN(n361) );
  XNOR2_X1 U350 ( .A(n263), .B(a[6]), .ZN(n254) );
  NOR2_X1 U351 ( .A1(n64), .A2(n61), .ZN(n3) );
  XOR2_X1 U352 ( .A(n74), .B(n363), .Z(product[7]) );
  NAND2_X1 U353 ( .A1(n105), .A2(n73), .ZN(n363) );
  XNOR2_X1 U354 ( .A(n264), .B(a[4]), .ZN(n255) );
  INV_X1 U355 ( .A(n30), .ZN(n28) );
  XNOR2_X1 U356 ( .A(n370), .B(n364), .ZN(product[9]) );
  AND2_X1 U357 ( .A1(n103), .A2(n65), .ZN(n364) );
  INV_X1 U358 ( .A(n31), .ZN(n29) );
  NAND2_X1 U359 ( .A1(n52), .A2(n32), .ZN(n30) );
  INV_X1 U360 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U361 ( .A1(n309), .A2(n21), .ZN(n19) );
  NAND2_X1 U362 ( .A1(n309), .A2(n39), .ZN(n37) );
  NAND2_X1 U363 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U364 ( .A1(n309), .A2(n28), .ZN(n26) );
  INV_X1 U365 ( .A(n3), .ZN(n57) );
  NAND2_X1 U366 ( .A1(n100), .A2(n44), .ZN(n6) );
  XNOR2_X1 U367 ( .A(n321), .B(n13), .ZN(product[5]) );
  NAND2_X1 U368 ( .A1(n319), .A2(n82), .ZN(n13) );
  XNOR2_X1 U369 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U370 ( .A1(n365), .A2(n94), .ZN(n16) );
  NOR2_X1 U371 ( .A1(n41), .A2(n34), .ZN(n32) );
  NAND2_X1 U372 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U373 ( .A(n61), .ZN(n102) );
  XNOR2_X1 U374 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U375 ( .A1(n52), .A2(n51), .ZN(n7) );
  AOI21_X1 U376 ( .B1(n365), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U377 ( .A(n94), .ZN(n92) );
  XNOR2_X1 U378 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U379 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U380 ( .A(n34), .ZN(n99) );
  NOR2_X1 U381 ( .A1(n50), .A2(n41), .ZN(n39) );
  INV_X1 U382 ( .A(n50), .ZN(n52) );
  NAND2_X1 U383 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U384 ( .A(n349), .ZN(n104) );
  AOI21_X1 U385 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U386 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  AOI21_X1 U387 ( .B1(n366), .B2(n83), .A(n334), .ZN(n78) );
  NOR2_X1 U388 ( .A1(n125), .A2(n130), .ZN(n64) );
  XOR2_X1 U389 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U390 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U391 ( .A(n84), .ZN(n108) );
  OAI21_X1 U392 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  NAND2_X1 U393 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U394 ( .A(n23), .ZN(n98) );
  OAI21_X1 U395 ( .B1(n311), .B2(n76), .A(n77), .ZN(n75) );
  NOR2_X1 U396 ( .A1(n30), .A2(n23), .ZN(n21) );
  NAND2_X1 U397 ( .A1(n125), .A2(n130), .ZN(n65) );
  XOR2_X1 U398 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U399 ( .A(n88), .ZN(n109) );
  OAI21_X1 U400 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U401 ( .A(n51), .ZN(n53) );
  NAND2_X1 U402 ( .A1(n131), .A2(n136), .ZN(n70) );
  XOR2_X1 U403 ( .A(n12), .B(n328), .Z(product[6]) );
  NAND2_X1 U404 ( .A1(n346), .A2(n77), .ZN(n12) );
  XNOR2_X1 U405 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U406 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U407 ( .A1(n116), .A2(n115), .ZN(n41) );
  NOR2_X1 U408 ( .A1(n170), .A2(n112), .ZN(n23) );
  INV_X1 U409 ( .A(n112), .ZN(n113) );
  NOR2_X1 U410 ( .A1(n114), .A2(n113), .ZN(n34) );
  OR2_X1 U411 ( .A1(n200), .A2(n193), .ZN(n365) );
  NAND2_X1 U412 ( .A1(n170), .A2(n112), .ZN(n24) );
  NOR2_X1 U413 ( .A1(n137), .A2(n142), .ZN(n72) );
  NOR2_X1 U414 ( .A1(n117), .A2(n120), .ZN(n50) );
  NOR2_X1 U415 ( .A1(n151), .A2(n331), .ZN(n84) );
  NOR2_X1 U416 ( .A1(n143), .A2(n146), .ZN(n76) );
  OR2_X1 U417 ( .A1(n147), .A2(n150), .ZN(n366) );
  NAND2_X1 U418 ( .A1(n116), .A2(n115), .ZN(n44) );
  NAND2_X1 U419 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U420 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U421 ( .A1(n117), .A2(n120), .ZN(n51) );
  INV_X1 U422 ( .A(n97), .ZN(n95) );
  NAND2_X1 U423 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U424 ( .A1(n147), .A2(n150), .ZN(n82) );
  NAND2_X1 U425 ( .A1(n143), .A2(n146), .ZN(n77) );
  NAND2_X1 U426 ( .A1(n151), .A2(n331), .ZN(n85) );
  AND2_X1 U427 ( .A1(n323), .A2(n161), .ZN(n193) );
  OR2_X1 U428 ( .A1(n374), .A2(n260), .ZN(n228) );
  OR2_X1 U429 ( .A1(n374), .A2(n259), .ZN(n219) );
  OAI22_X1 U430 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  INV_X1 U431 ( .A(n118), .ZN(n119) );
  OAI22_X1 U432 ( .A1(n307), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  AND2_X1 U433 ( .A1(n374), .A2(n158), .ZN(n185) );
  OAI22_X1 U434 ( .A1(n308), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  INV_X1 U435 ( .A(n157), .ZN(n178) );
  INV_X1 U436 ( .A(n163), .ZN(n194) );
  OAI22_X1 U437 ( .A1(n229), .A2(n308), .B1(n229), .B2(n273), .ZN(n163) );
  OAI22_X1 U438 ( .A1(n307), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  AND2_X1 U439 ( .A1(n323), .A2(n155), .ZN(n177) );
  OAI22_X1 U440 ( .A1(n308), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  INV_X1 U441 ( .A(n154), .ZN(n170) );
  OR2_X1 U442 ( .A1(n323), .A2(n258), .ZN(n210) );
  AND2_X1 U443 ( .A1(n332), .A2(n97), .ZN(product[1]) );
  OAI22_X1 U444 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OAI22_X1 U445 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OR2_X1 U446 ( .A1(n374), .A2(n261), .ZN(n237) );
  NAND2_X1 U447 ( .A1(n246), .A2(n254), .ZN(n250) );
  NAND2_X1 U448 ( .A1(n310), .A2(n248), .ZN(n252) );
  AND2_X1 U449 ( .A1(n323), .A2(n164), .ZN(product[0]) );
  BUF_X2 U450 ( .A(n1), .Z(n370) );
  AOI21_X1 U451 ( .B1(n67), .B2(n312), .A(n68), .ZN(n1) );
  NAND2_X1 U452 ( .A1(n200), .A2(n193), .ZN(n94) );
  OAI22_X1 U453 ( .A1(n307), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  XNOR2_X1 U454 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U455 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U456 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U457 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U458 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U459 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U460 ( .A(n262), .B(n374), .ZN(n209) );
  INV_X1 U461 ( .A(n262), .ZN(n258) );
  XNOR2_X1 U462 ( .A(b[1]), .B(n262), .ZN(n208) );
  XNOR2_X1 U463 ( .A(n265), .B(a[2]), .ZN(n256) );
  XNOR2_X1 U464 ( .A(n63), .B(n8), .ZN(product[10]) );
  INV_X1 U465 ( .A(n87), .ZN(n86) );
  NOR2_X1 U466 ( .A1(n153), .A2(n168), .ZN(n88) );
  NOR2_X1 U467 ( .A1(n72), .A2(n349), .ZN(n67) );
  XNOR2_X1 U468 ( .A(n71), .B(n10), .ZN(product[8]) );
  OAI21_X1 U469 ( .B1(n320), .B2(n72), .A(n304), .ZN(n71) );
  AOI21_X1 U470 ( .B1(n325), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U471 ( .B1(n325), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U472 ( .A(n325), .ZN(n58) );
  AOI21_X1 U473 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U474 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  INV_X1 U475 ( .A(n128), .ZN(n129) );
  INV_X1 U476 ( .A(n160), .ZN(n186) );
  OAI21_X1 U477 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  INV_X1 U478 ( .A(n41), .ZN(n100) );
  OAI21_X1 U479 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NAND2_X1 U480 ( .A1(n109), .A2(n89), .ZN(n15) );
  NAND2_X1 U481 ( .A1(n153), .A2(n168), .ZN(n89) );
  INV_X1 U482 ( .A(n312), .ZN(n74) );
  NAND2_X1 U483 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI21_X1 U484 ( .B1(n370), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U485 ( .B1(n370), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U486 ( .B1(n369), .B2(n64), .A(n65), .ZN(n63) );
  OAI21_X1 U487 ( .B1(n370), .B2(n57), .A(n58), .ZN(n56) );
  OAI22_X1 U488 ( .A1(n202), .A2(n361), .B1(n202), .B2(n351), .ZN(n154) );
  OAI22_X1 U489 ( .A1(n361), .A2(n206), .B1(n205), .B2(n351), .ZN(n173) );
  OAI22_X1 U490 ( .A1(n360), .A2(n203), .B1(n202), .B2(n351), .ZN(n112) );
  OAI22_X1 U491 ( .A1(n361), .A2(n205), .B1(n204), .B2(n351), .ZN(n172) );
  OAI22_X1 U492 ( .A1(n360), .A2(n204), .B1(n203), .B2(n351), .ZN(n171) );
  OAI22_X1 U493 ( .A1(n360), .A2(n207), .B1(n206), .B2(n351), .ZN(n174) );
  OAI22_X1 U494 ( .A1(n361), .A2(n208), .B1(n207), .B2(n351), .ZN(n175) );
  INV_X1 U495 ( .A(n362), .ZN(n155) );
  XNOR2_X1 U496 ( .A(b[5]), .B(n345), .ZN(n213) );
  OAI22_X1 U497 ( .A1(n250), .A2(n258), .B1(n210), .B2(n362), .ZN(n166) );
  OAI22_X1 U498 ( .A1(n250), .A2(n209), .B1(n208), .B2(n362), .ZN(n176) );
  XNOR2_X1 U499 ( .A(b[6]), .B(n322), .ZN(n212) );
  XNOR2_X1 U500 ( .A(b[7]), .B(n345), .ZN(n211) );
  XNOR2_X1 U501 ( .A(b[4]), .B(n322), .ZN(n214) );
  XNOR2_X1 U502 ( .A(b[2]), .B(n303), .ZN(n216) );
  XNOR2_X1 U503 ( .A(b[3]), .B(n303), .ZN(n215) );
  XNOR2_X1 U504 ( .A(n303), .B(n323), .ZN(n218) );
  XNOR2_X1 U505 ( .A(b[1]), .B(n263), .ZN(n217) );
  INV_X1 U506 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U507 ( .A(n25), .B(n4), .ZN(product[14]) );
  OAI21_X1 U508 ( .B1(n370), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U509 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  XNOR2_X1 U510 ( .A(n45), .B(n6), .ZN(product[12]) );
  OAI21_X1 U511 ( .B1(n370), .B2(n46), .A(n47), .ZN(n45) );
  OAI22_X1 U512 ( .A1(n352), .A2(n217), .B1(n216), .B2(n372), .ZN(n183) );
  OAI22_X1 U513 ( .A1(n353), .A2(n212), .B1(n211), .B2(n306), .ZN(n118) );
  OAI22_X1 U514 ( .A1(n211), .A2(n352), .B1(n211), .B2(n306), .ZN(n157) );
  OAI22_X1 U515 ( .A1(n352), .A2(n213), .B1(n212), .B2(n372), .ZN(n179) );
  OAI22_X1 U516 ( .A1(n353), .A2(n214), .B1(n213), .B2(n372), .ZN(n180) );
  OAI22_X1 U517 ( .A1(n353), .A2(n216), .B1(n215), .B2(n372), .ZN(n182) );
  OAI22_X1 U518 ( .A1(n352), .A2(n215), .B1(n214), .B2(n372), .ZN(n181) );
  INV_X1 U519 ( .A(n372), .ZN(n158) );
  XNOR2_X1 U520 ( .A(b[4]), .B(n348), .ZN(n223) );
  XNOR2_X1 U521 ( .A(n348), .B(b[5]), .ZN(n222) );
  XNOR2_X1 U522 ( .A(n348), .B(b[6]), .ZN(n221) );
  OAI22_X1 U523 ( .A1(n251), .A2(n259), .B1(n219), .B2(n372), .ZN(n167) );
  XNOR2_X1 U524 ( .A(b[3]), .B(n348), .ZN(n224) );
  OAI22_X1 U525 ( .A1(n251), .A2(n218), .B1(n217), .B2(n372), .ZN(n184) );
  XNOR2_X1 U526 ( .A(b[7]), .B(n347), .ZN(n220) );
  INV_X1 U527 ( .A(n348), .ZN(n260) );
  XNOR2_X1 U528 ( .A(b[2]), .B(n348), .ZN(n225) );
  XNOR2_X1 U529 ( .A(n348), .B(n323), .ZN(n227) );
  XNOR2_X1 U530 ( .A(b[1]), .B(n347), .ZN(n226) );
  OAI22_X1 U531 ( .A1(n339), .A2(n221), .B1(n220), .B2(n373), .ZN(n128) );
  OAI22_X1 U532 ( .A1(n220), .A2(n358), .B1(n220), .B2(n326), .ZN(n160) );
  OAI22_X1 U533 ( .A1(n359), .A2(n305), .B1(n221), .B2(n326), .ZN(n187) );
  OAI22_X1 U534 ( .A1(n223), .A2(n359), .B1(n222), .B2(n373), .ZN(n188) );
  OAI22_X1 U535 ( .A1(n358), .A2(n225), .B1(n224), .B2(n326), .ZN(n190) );
  OAI22_X1 U536 ( .A1(n358), .A2(n224), .B1(n326), .B2(n223), .ZN(n189) );
  OAI22_X1 U537 ( .A1(n339), .A2(n226), .B1(n225), .B2(n373), .ZN(n191) );
  OAI22_X1 U538 ( .A1(n359), .A2(n260), .B1(n228), .B2(n373), .ZN(n168) );
  XNOR2_X1 U539 ( .A(n330), .B(b[5]), .ZN(n231) );
  XNOR2_X1 U540 ( .A(b[6]), .B(n265), .ZN(n230) );
  XNOR2_X1 U541 ( .A(n318), .B(b[4]), .ZN(n232) );
  INV_X1 U542 ( .A(n350), .ZN(n161) );
  OAI22_X1 U543 ( .A1(n252), .A2(n227), .B1(n256), .B2(n226), .ZN(n192) );
  XNOR2_X1 U544 ( .A(b[7]), .B(n265), .ZN(n229) );
  XNOR2_X1 U545 ( .A(n318), .B(n374), .ZN(n236) );
  XNOR2_X1 U546 ( .A(b[2]), .B(n265), .ZN(n234) );
  XNOR2_X1 U547 ( .A(b[3]), .B(n265), .ZN(n233) );
  INV_X1 U548 ( .A(n265), .ZN(n261) );
  XNOR2_X1 U549 ( .A(b[1]), .B(n265), .ZN(n235) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n80, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102, n103,
         n105, n106, n108, n109, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n157, n158, n160, n161, n163, n164, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n245, n246, n248, n249, n250, n251, n252,
         n253, n255, n256, n258, n259, n260, n261, n262, n263, n264, n265,
         n273, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n360, n361, n362;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U141 ( .A(n195), .B(n188), .CI(n182), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  CLKBUF_X1 U268 ( .A(n265), .Z(n303) );
  CLKBUF_X1 U269 ( .A(n141), .Z(n304) );
  CLKBUF_X1 U270 ( .A(n265), .Z(n305) );
  BUF_X1 U271 ( .A(n333), .Z(n306) );
  CLKBUF_X1 U272 ( .A(n265), .Z(n307) );
  CLKBUF_X1 U273 ( .A(n265), .Z(n308) );
  XNOR2_X1 U274 ( .A(n265), .B(n334), .ZN(n309) );
  XOR2_X1 U275 ( .A(n141), .B(n144), .Z(n310) );
  XOR2_X1 U276 ( .A(n139), .B(n310), .Z(n137) );
  NAND2_X1 U277 ( .A1(n139), .A2(n304), .ZN(n311) );
  NAND2_X1 U278 ( .A1(n139), .A2(n144), .ZN(n312) );
  NAND2_X1 U279 ( .A1(n141), .A2(n144), .ZN(n313) );
  NAND3_X1 U280 ( .A1(n311), .A2(n312), .A3(n313), .ZN(n136) );
  CLKBUF_X1 U281 ( .A(n90), .Z(n314) );
  OAI21_X1 U282 ( .B1(n84), .B2(n86), .A(n85), .ZN(n315) );
  NAND2_X1 U283 ( .A1(n317), .A2(n146), .ZN(n316) );
  FA_X1 U284 ( .A(n148), .B(n183), .CI(n145), .S(n317) );
  CLKBUF_X1 U285 ( .A(n263), .Z(n318) );
  OAI22_X1 U286 ( .A1(n335), .A2(n261), .B1(n237), .B2(n273), .ZN(n319) );
  XOR2_X1 U287 ( .A(n184), .B(n167), .Z(n320) );
  NAND2_X1 U288 ( .A1(n249), .A2(n273), .ZN(n321) );
  CLKBUF_X1 U289 ( .A(n265), .Z(n338) );
  BUF_X2 U290 ( .A(n264), .Z(n322) );
  BUF_X1 U291 ( .A(n133), .Z(n323) );
  OAI21_X1 U292 ( .B1(n347), .B2(n73), .A(n70), .ZN(n324) );
  XOR2_X1 U293 ( .A(n263), .B(a[6]), .Z(n325) );
  XOR2_X1 U294 ( .A(n190), .B(n197), .Z(n326) );
  XOR2_X1 U295 ( .A(n149), .B(n326), .Z(n147) );
  NAND2_X1 U296 ( .A1(n320), .A2(n190), .ZN(n327) );
  NAND2_X1 U297 ( .A1(n320), .A2(n197), .ZN(n328) );
  NAND2_X1 U298 ( .A1(n190), .A2(n197), .ZN(n329) );
  NAND3_X1 U299 ( .A1(n327), .A2(n328), .A3(n329), .ZN(n146) );
  BUF_X2 U300 ( .A(n340), .Z(n330) );
  NOR2_X2 U301 ( .A1(n121), .A2(n124), .ZN(n61) );
  OR2_X1 U302 ( .A1(n131), .A2(n136), .ZN(n331) );
  OR2_X1 U303 ( .A1(n201), .A2(n319), .ZN(n332) );
  BUF_X2 U304 ( .A(n256), .Z(n360) );
  XNOR2_X1 U305 ( .A(n263), .B(a[6]), .ZN(n333) );
  INV_X1 U306 ( .A(n164), .ZN(n334) );
  NAND2_X1 U307 ( .A1(n309), .A2(n273), .ZN(n335) );
  NAND2_X1 U308 ( .A1(n249), .A2(n273), .ZN(n253) );
  INV_X1 U309 ( .A(n103), .ZN(n336) );
  NAND2_X1 U310 ( .A1(n246), .A2(n333), .ZN(n337) );
  XNOR2_X1 U311 ( .A(n133), .B(n339), .ZN(n131) );
  XNOR2_X1 U312 ( .A(n135), .B(n138), .ZN(n339) );
  XNOR2_X1 U313 ( .A(n264), .B(a[4]), .ZN(n340) );
  INV_X1 U314 ( .A(n260), .ZN(n341) );
  NAND2_X1 U315 ( .A1(n323), .A2(n135), .ZN(n342) );
  NAND2_X1 U316 ( .A1(n323), .A2(n138), .ZN(n343) );
  NAND2_X1 U317 ( .A1(n135), .A2(n138), .ZN(n344) );
  NAND3_X1 U318 ( .A1(n342), .A2(n343), .A3(n344), .ZN(n130) );
  XNOR2_X1 U319 ( .A(n265), .B(n334), .ZN(n249) );
  OAI21_X1 U320 ( .B1(n61), .B2(n65), .A(n62), .ZN(n345) );
  OAI21_X1 U321 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  XNOR2_X1 U322 ( .A(n265), .B(a[2]), .ZN(n346) );
  NOR2_X1 U323 ( .A1(n131), .A2(n136), .ZN(n347) );
  NOR2_X1 U324 ( .A1(n131), .A2(n136), .ZN(n348) );
  CLKBUF_X1 U325 ( .A(n256), .Z(n361) );
  NOR2_X2 U326 ( .A1(n64), .A2(n61), .ZN(n3) );
  NOR2_X1 U327 ( .A1(n317), .A2(n146), .ZN(n349) );
  INV_X1 U328 ( .A(n325), .ZN(n350) );
  NOR2_X1 U329 ( .A1(n143), .A2(n146), .ZN(n76) );
  AOI21_X1 U330 ( .B1(n315), .B2(n358), .A(n80), .ZN(n351) );
  NAND2_X1 U331 ( .A1(n356), .A2(n255), .ZN(n352) );
  OAI21_X1 U332 ( .B1(n349), .B2(n351), .A(n316), .ZN(n353) );
  NAND2_X1 U333 ( .A1(n248), .A2(n346), .ZN(n354) );
  AOI21_X2 U334 ( .B1(n67), .B2(n353), .A(n324), .ZN(n355) );
  AOI21_X1 U335 ( .B1(n67), .B2(n353), .A(n324), .ZN(n1) );
  BUF_X2 U336 ( .A(n245), .Z(n362) );
  INV_X2 U337 ( .A(n164), .ZN(n273) );
  NAND2_X1 U338 ( .A1(n356), .A2(n255), .ZN(n251) );
  XOR2_X1 U339 ( .A(n263), .B(a[4]), .Z(n356) );
  INV_X1 U340 ( .A(n30), .ZN(n28) );
  NAND2_X1 U341 ( .A1(n103), .A2(n65), .ZN(n9) );
  INV_X1 U342 ( .A(n64), .ZN(n103) );
  INV_X1 U343 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U344 ( .A1(n3), .A2(n21), .ZN(n19) );
  INV_X1 U345 ( .A(n31), .ZN(n29) );
  NAND2_X1 U346 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U347 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U348 ( .A1(n3), .A2(n28), .ZN(n26) );
  NAND2_X1 U349 ( .A1(n3), .A2(n39), .ZN(n37) );
  INV_X1 U350 ( .A(n3), .ZN(n57) );
  NAND2_X1 U351 ( .A1(n52), .A2(n51), .ZN(n7) );
  XNOR2_X1 U352 ( .A(n13), .B(n315), .ZN(product[5]) );
  NAND2_X1 U353 ( .A1(n358), .A2(n82), .ZN(n13) );
  XNOR2_X1 U354 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U355 ( .A1(n357), .A2(n94), .ZN(n16) );
  NAND2_X1 U356 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U357 ( .A(n61), .ZN(n102) );
  XNOR2_X1 U358 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U359 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U360 ( .A(n23), .ZN(n98) );
  AOI21_X1 U361 ( .B1(n83), .B2(n358), .A(n80), .ZN(n78) );
  INV_X1 U362 ( .A(n82), .ZN(n80) );
  NAND2_X1 U363 ( .A1(n105), .A2(n73), .ZN(n11) );
  INV_X1 U364 ( .A(n72), .ZN(n105) );
  XNOR2_X1 U365 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U366 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U367 ( .A(n41), .ZN(n100) );
  XNOR2_X1 U368 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U369 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U370 ( .A(n34), .ZN(n99) );
  AOI21_X1 U371 ( .B1(n357), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U372 ( .A(n94), .ZN(n92) );
  INV_X1 U373 ( .A(n50), .ZN(n52) );
  NAND2_X1 U374 ( .A1(n331), .A2(n70), .ZN(n10) );
  AOI21_X1 U375 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U376 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  OAI21_X1 U377 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  NOR2_X1 U378 ( .A1(n125), .A2(n130), .ZN(n64) );
  NOR2_X1 U379 ( .A1(n41), .A2(n34), .ZN(n32) );
  OAI21_X1 U380 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  NOR2_X1 U381 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U382 ( .A1(n50), .A2(n41), .ZN(n39) );
  NAND2_X1 U383 ( .A1(n125), .A2(n130), .ZN(n65) );
  OAI21_X1 U384 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U385 ( .A(n51), .ZN(n53) );
  NAND2_X1 U386 ( .A1(n131), .A2(n136), .ZN(n70) );
  XOR2_X1 U387 ( .A(n12), .B(n351), .Z(product[6]) );
  NAND2_X1 U388 ( .A1(n106), .A2(n316), .ZN(n12) );
  INV_X1 U389 ( .A(n349), .ZN(n106) );
  XOR2_X1 U390 ( .A(n15), .B(n314), .Z(product[3]) );
  NAND2_X1 U391 ( .A1(n109), .A2(n89), .ZN(n15) );
  INV_X1 U392 ( .A(n88), .ZN(n109) );
  NOR2_X1 U393 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U394 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U395 ( .A1(n187), .A2(n175), .ZN(n134) );
  OAI21_X1 U396 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  NOR2_X1 U397 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U398 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U399 ( .A(n112), .ZN(n113) );
  XOR2_X1 U400 ( .A(n14), .B(n86), .Z(product[4]) );
  INV_X1 U401 ( .A(n84), .ZN(n108) );
  NOR2_X1 U402 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U403 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U404 ( .A1(n116), .A2(n115), .ZN(n44) );
  INV_X1 U405 ( .A(n97), .ZN(n95) );
  NOR2_X1 U406 ( .A1(n137), .A2(n142), .ZN(n72) );
  OR2_X1 U407 ( .A1(n200), .A2(n193), .ZN(n357) );
  NAND2_X1 U408 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U409 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U410 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U411 ( .A1(n147), .A2(n150), .ZN(n82) );
  NAND2_X1 U412 ( .A1(n143), .A2(n146), .ZN(n77) );
  OR2_X1 U413 ( .A1(n150), .A2(n147), .ZN(n358) );
  OAI21_X1 U414 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NAND2_X1 U415 ( .A1(n121), .A2(n124), .ZN(n62) );
  AND2_X1 U416 ( .A1(n362), .A2(n161), .ZN(n193) );
  AND2_X1 U417 ( .A1(n362), .A2(n158), .ZN(n185) );
  INV_X1 U418 ( .A(n157), .ZN(n178) );
  INV_X1 U419 ( .A(n118), .ZN(n119) );
  NOR2_X1 U420 ( .A1(n153), .A2(n168), .ZN(n88) );
  OR2_X1 U421 ( .A1(n362), .A2(n259), .ZN(n219) );
  AND2_X1 U422 ( .A1(n332), .A2(n97), .ZN(product[1]) );
  NOR2_X1 U423 ( .A1(n151), .A2(n152), .ZN(n84) );
  INV_X1 U424 ( .A(n128), .ZN(n129) );
  INV_X1 U425 ( .A(n163), .ZN(n194) );
  INV_X1 U426 ( .A(n160), .ZN(n186) );
  AND2_X1 U427 ( .A1(n362), .A2(n325), .ZN(n177) );
  INV_X1 U428 ( .A(n154), .ZN(n170) );
  OR2_X1 U429 ( .A1(n362), .A2(n258), .ZN(n210) );
  NAND2_X1 U430 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U431 ( .A1(n362), .A2(n260), .ZN(n228) );
  OR2_X1 U432 ( .A1(n362), .A2(n261), .ZN(n237) );
  NAND2_X1 U433 ( .A1(n248), .A2(n346), .ZN(n252) );
  NAND2_X1 U434 ( .A1(n246), .A2(n333), .ZN(n250) );
  AND2_X1 U435 ( .A1(n362), .A2(n164), .ZN(product[0]) );
  OAI22_X1 U436 ( .A1(n335), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  OAI22_X1 U437 ( .A1(n335), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  OAI22_X1 U438 ( .A1(n321), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U439 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U440 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U441 ( .A1(n321), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OAI22_X1 U442 ( .A1(n229), .A2(n335), .B1(n229), .B2(n273), .ZN(n163) );
  OAI22_X1 U443 ( .A1(n321), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  NOR2_X1 U444 ( .A1(n348), .A2(n72), .ZN(n67) );
  XNOR2_X1 U445 ( .A(b[3]), .B(n263), .ZN(n215) );
  XNOR2_X1 U446 ( .A(b[7]), .B(n318), .ZN(n211) );
  XNOR2_X1 U447 ( .A(b[4]), .B(n318), .ZN(n214) );
  XNOR2_X1 U448 ( .A(b[5]), .B(n263), .ZN(n213) );
  AOI21_X1 U449 ( .B1(n345), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U450 ( .B1(n345), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U451 ( .B1(n345), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U452 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  INV_X1 U453 ( .A(n2), .ZN(n58) );
  XNOR2_X1 U454 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U455 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U456 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U457 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U458 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U459 ( .A(n262), .B(n362), .ZN(n209) );
  INV_X1 U460 ( .A(n262), .ZN(n258) );
  XOR2_X1 U461 ( .A(a[6]), .B(n262), .Z(n246) );
  XNOR2_X1 U462 ( .A(n264), .B(a[4]), .ZN(n255) );
  XNOR2_X1 U463 ( .A(n265), .B(a[2]), .ZN(n256) );
  XNOR2_X1 U464 ( .A(n63), .B(n8), .ZN(product[10]) );
  XNOR2_X1 U465 ( .A(n71), .B(n10), .ZN(product[8]) );
  XNOR2_X1 U466 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U467 ( .A1(n200), .A2(n193), .ZN(n94) );
  XNOR2_X1 U468 ( .A(b[2]), .B(n263), .ZN(n216) );
  XNOR2_X1 U469 ( .A(b[2]), .B(n262), .ZN(n207) );
  NAND2_X1 U470 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U471 ( .A1(n335), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  XNOR2_X1 U472 ( .A(b[1]), .B(n262), .ZN(n208) );
  NAND2_X1 U473 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U474 ( .A(n87), .ZN(n86) );
  INV_X1 U475 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U476 ( .A(b[1]), .B(n263), .ZN(n217) );
  XNOR2_X1 U477 ( .A(n263), .B(n362), .ZN(n218) );
  XNOR2_X1 U478 ( .A(b[6]), .B(n263), .ZN(n212) );
  XOR2_X1 U479 ( .A(n74), .B(n11), .Z(product[7]) );
  OAI21_X1 U480 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  OAI22_X1 U481 ( .A1(n252), .A2(n222), .B1(n221), .B2(n360), .ZN(n187) );
  OAI22_X1 U482 ( .A1(n252), .A2(n223), .B1(n222), .B2(n360), .ZN(n188) );
  OAI22_X1 U483 ( .A1(n252), .A2(n225), .B1(n224), .B2(n361), .ZN(n190) );
  OAI22_X1 U484 ( .A1(n252), .A2(n260), .B1(n228), .B2(n360), .ZN(n168) );
  OAI22_X1 U485 ( .A1(n354), .A2(n221), .B1(n220), .B2(n360), .ZN(n128) );
  OAI22_X1 U486 ( .A1(n354), .A2(n224), .B1(n223), .B2(n360), .ZN(n189) );
  OAI22_X1 U487 ( .A1(n220), .A2(n252), .B1(n220), .B2(n361), .ZN(n160) );
  OAI22_X1 U488 ( .A1(n252), .A2(n226), .B1(n225), .B2(n361), .ZN(n191) );
  OAI22_X1 U489 ( .A1(n354), .A2(n227), .B1(n226), .B2(n360), .ZN(n192) );
  XNOR2_X1 U490 ( .A(b[7]), .B(n338), .ZN(n229) );
  XNOR2_X1 U491 ( .A(b[5]), .B(n303), .ZN(n231) );
  INV_X1 U492 ( .A(n361), .ZN(n161) );
  XNOR2_X1 U493 ( .A(b[6]), .B(n265), .ZN(n230) );
  XNOR2_X1 U494 ( .A(b[4]), .B(n338), .ZN(n232) );
  XNOR2_X1 U495 ( .A(b[3]), .B(n307), .ZN(n233) );
  XNOR2_X1 U496 ( .A(n308), .B(n362), .ZN(n236) );
  XNOR2_X1 U497 ( .A(b[2]), .B(n338), .ZN(n234) );
  XNOR2_X1 U498 ( .A(b[1]), .B(n307), .ZN(n235) );
  INV_X1 U499 ( .A(n305), .ZN(n261) );
  OAI21_X1 U500 ( .B1(n355), .B2(n19), .A(n20), .ZN(n18) );
  XOR2_X1 U501 ( .A(n1), .B(n9), .Z(product[9]) );
  OAI21_X1 U502 ( .B1(n355), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U503 ( .B1(n355), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U504 ( .B1(n355), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U505 ( .B1(n355), .B2(n26), .A(n27), .ZN(n25) );
  OAI22_X1 U506 ( .A1(n202), .A2(n337), .B1(n202), .B2(n350), .ZN(n154) );
  OAI22_X1 U507 ( .A1(n337), .A2(n206), .B1(n205), .B2(n350), .ZN(n173) );
  OAI22_X1 U508 ( .A1(n337), .A2(n203), .B1(n202), .B2(n350), .ZN(n112) );
  OAI22_X1 U509 ( .A1(n337), .A2(n205), .B1(n204), .B2(n350), .ZN(n172) );
  OAI22_X1 U510 ( .A1(n337), .A2(n208), .B1(n207), .B2(n350), .ZN(n175) );
  OAI22_X1 U511 ( .A1(n337), .A2(n204), .B1(n203), .B2(n350), .ZN(n171) );
  OAI22_X1 U512 ( .A1(n337), .A2(n207), .B1(n206), .B2(n306), .ZN(n174) );
  OAI22_X1 U513 ( .A1(n250), .A2(n258), .B1(n210), .B2(n306), .ZN(n166) );
  OAI22_X1 U514 ( .A1(n250), .A2(n209), .B1(n208), .B2(n306), .ZN(n176) );
  OAI22_X1 U515 ( .A1(n251), .A2(n217), .B1(n216), .B2(n330), .ZN(n183) );
  OAI22_X1 U516 ( .A1(n251), .A2(n215), .B1(n214), .B2(n330), .ZN(n181) );
  OAI22_X1 U517 ( .A1(n352), .A2(n212), .B1(n211), .B2(n330), .ZN(n118) );
  OAI22_X1 U518 ( .A1(n251), .A2(n216), .B1(n215), .B2(n340), .ZN(n182) );
  OAI22_X1 U519 ( .A1(n251), .A2(n214), .B1(n213), .B2(n330), .ZN(n180) );
  OAI22_X1 U520 ( .A1(n211), .A2(n352), .B1(n211), .B2(n330), .ZN(n157) );
  OAI22_X1 U521 ( .A1(n251), .A2(n213), .B1(n212), .B2(n340), .ZN(n179) );
  INV_X1 U522 ( .A(n340), .ZN(n158) );
  OAI22_X1 U523 ( .A1(n352), .A2(n259), .B1(n219), .B2(n340), .ZN(n167) );
  OAI22_X1 U524 ( .A1(n352), .A2(n218), .B1(n217), .B2(n340), .ZN(n184) );
  INV_X1 U525 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U526 ( .A(b[5]), .B(n341), .ZN(n222) );
  XNOR2_X1 U527 ( .A(b[3]), .B(n322), .ZN(n224) );
  XNOR2_X1 U528 ( .A(b[4]), .B(n322), .ZN(n223) );
  XNOR2_X1 U529 ( .A(b[2]), .B(n322), .ZN(n225) );
  XNOR2_X1 U530 ( .A(b[6]), .B(n341), .ZN(n221) );
  XNOR2_X1 U531 ( .A(n322), .B(n362), .ZN(n227) );
  XNOR2_X1 U532 ( .A(b[1]), .B(n322), .ZN(n226) );
  XNOR2_X1 U533 ( .A(b[7]), .B(n322), .ZN(n220) );
  XOR2_X1 U534 ( .A(n264), .B(a[2]), .Z(n248) );
  INV_X1 U535 ( .A(n75), .ZN(n74) );
  NAND2_X1 U536 ( .A1(n153), .A2(n168), .ZN(n89) );
  OAI21_X1 U537 ( .B1(n1), .B2(n336), .A(n65), .ZN(n63) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n80, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n92, n94, n97, n98, n99, n100, n103, n105,
         n106, n108, n109, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n157, n158, n160, n161, n163, n164, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n245, n248, n249, n250, n252, n253, n255, n256,
         n258, n259, n260, n261, n262, n263, n264, n265, n273, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n361, n362, n363;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n186), .CI(n128), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n177), .B(n189), .CI(n196), .CO(n144), .S(n145) );
  HA_X1 U146 ( .A(n167), .B(n184), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n199), .B(n192), .CO(n152), .S(n153) );
  CLKBUF_X1 U268 ( .A(n264), .Z(n303) );
  OAI21_X1 U269 ( .B1(n84), .B2(n86), .A(n85), .ZN(n304) );
  CLKBUF_X1 U270 ( .A(n353), .Z(n305) );
  AND2_X2 U271 ( .A1(n201), .A2(n169), .ZN(n306) );
  INV_X4 U272 ( .A(n306), .ZN(n97) );
  XNOR2_X1 U273 ( .A(n133), .B(n307), .ZN(n131) );
  XNOR2_X1 U274 ( .A(n138), .B(n135), .ZN(n307) );
  NOR2_X1 U275 ( .A1(n64), .A2(n336), .ZN(n308) );
  CLKBUF_X1 U276 ( .A(n264), .Z(n309) );
  NOR2_X1 U277 ( .A1(n64), .A2(n336), .ZN(n3) );
  CLKBUF_X1 U278 ( .A(n121), .Z(n310) );
  BUF_X2 U279 ( .A(n362), .Z(n311) );
  BUF_X2 U280 ( .A(n256), .Z(n362) );
  CLKBUF_X1 U281 ( .A(b[3]), .Z(n318) );
  OR2_X1 U282 ( .A1(n310), .A2(n124), .ZN(n312) );
  CLKBUF_X1 U283 ( .A(n264), .Z(n313) );
  NAND2_X1 U284 ( .A1(n248), .A2(n361), .ZN(n353) );
  CLKBUF_X1 U285 ( .A(n86), .Z(n314) );
  CLKBUF_X1 U286 ( .A(n224), .Z(n315) );
  CLKBUF_X1 U287 ( .A(n89), .Z(n316) );
  XNOR2_X1 U288 ( .A(n149), .B(n317), .ZN(n147) );
  XNOR2_X1 U289 ( .A(n190), .B(n197), .ZN(n317) );
  XOR2_X1 U290 ( .A(b[3]), .B(n259), .Z(n215) );
  OAI21_X1 U291 ( .B1(n338), .B2(n73), .A(n70), .ZN(n319) );
  OAI21_X1 U292 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  BUF_X2 U293 ( .A(n245), .Z(n363) );
  NOR2_X2 U294 ( .A1(n125), .A2(n130), .ZN(n64) );
  NAND2_X1 U295 ( .A1(n133), .A2(n138), .ZN(n320) );
  NAND2_X1 U296 ( .A1(n133), .A2(n135), .ZN(n321) );
  NAND2_X1 U297 ( .A1(n138), .A2(n135), .ZN(n322) );
  NAND3_X1 U298 ( .A1(n320), .A2(n321), .A3(n322), .ZN(n130) );
  NAND2_X1 U299 ( .A1(n357), .A2(n255), .ZN(n323) );
  NAND2_X1 U300 ( .A1(n149), .A2(n190), .ZN(n324) );
  NAND2_X1 U301 ( .A1(n149), .A2(n197), .ZN(n325) );
  NAND2_X1 U302 ( .A1(n190), .A2(n197), .ZN(n326) );
  NAND3_X1 U303 ( .A1(n324), .A2(n325), .A3(n326), .ZN(n146) );
  INV_X1 U304 ( .A(n259), .ZN(n327) );
  CLKBUF_X1 U305 ( .A(n263), .Z(n328) );
  OR2_X1 U306 ( .A1(n363), .A2(n261), .ZN(n237) );
  NAND2_X1 U307 ( .A1(n137), .A2(n142), .ZN(n73) );
  NOR2_X1 U308 ( .A1(n143), .A2(n146), .ZN(n76) );
  BUF_X1 U309 ( .A(n265), .Z(n335) );
  OR2_X1 U310 ( .A1(n131), .A2(n136), .ZN(n329) );
  OR2_X1 U311 ( .A1(n201), .A2(n169), .ZN(n330) );
  XOR2_X1 U312 ( .A(n263), .B(a[4]), .Z(n331) );
  INV_X1 U313 ( .A(n260), .ZN(n332) );
  XOR2_X1 U314 ( .A(n264), .B(a[2]), .Z(n333) );
  BUF_X2 U315 ( .A(n265), .Z(n334) );
  NOR2_X1 U316 ( .A1(n121), .A2(n124), .ZN(n336) );
  OAI21_X1 U317 ( .B1(n61), .B2(n65), .A(n62), .ZN(n337) );
  NOR2_X1 U318 ( .A1(n131), .A2(n136), .ZN(n338) );
  OR2_X2 U319 ( .A1(n343), .A2(n344), .ZN(n339) );
  NOR2_X1 U320 ( .A1(n131), .A2(n136), .ZN(n69) );
  OR2_X1 U321 ( .A1(n343), .A2(n344), .ZN(n250) );
  NOR2_X1 U322 ( .A1(n121), .A2(n124), .ZN(n61) );
  NAND2_X1 U323 ( .A1(n106), .A2(n77), .ZN(n12) );
  CLKBUF_X1 U324 ( .A(n263), .Z(n340) );
  NAND2_X1 U325 ( .A1(n331), .A2(n255), .ZN(n341) );
  NAND2_X1 U326 ( .A1(n331), .A2(n255), .ZN(n342) );
  OAI22_X1 U327 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OAI22_X1 U328 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  XNOR2_X2 U329 ( .A(n264), .B(a[4]), .ZN(n347) );
  INV_X1 U330 ( .A(n76), .ZN(n106) );
  XOR2_X1 U331 ( .A(n263), .B(a[6]), .Z(n343) );
  XNOR2_X1 U332 ( .A(a[6]), .B(n262), .ZN(n344) );
  AOI21_X1 U333 ( .B1(n356), .B2(n83), .A(n80), .ZN(n345) );
  AOI21_X1 U334 ( .B1(n304), .B2(n356), .A(n80), .ZN(n346) );
  XNOR2_X1 U335 ( .A(n354), .B(n348), .ZN(product[9]) );
  AND2_X1 U336 ( .A1(n103), .A2(n65), .ZN(n348) );
  BUF_X2 U337 ( .A(n355), .Z(n349) );
  BUF_X1 U338 ( .A(n355), .Z(n350) );
  AOI21_X1 U339 ( .B1(n67), .B2(n352), .A(n319), .ZN(n351) );
  AOI21_X1 U340 ( .B1(n67), .B2(n352), .A(n319), .ZN(n354) );
  OAI21_X1 U341 ( .B1(n346), .B2(n76), .A(n77), .ZN(n352) );
  AOI21_X1 U342 ( .B1(n67), .B2(n352), .A(n68), .ZN(n1) );
  XNOR2_X1 U343 ( .A(n263), .B(a[6]), .ZN(n355) );
  NOR2_X1 U344 ( .A1(n137), .A2(n142), .ZN(n72) );
  OR2_X1 U345 ( .A1(n147), .A2(n150), .ZN(n356) );
  OR2_X1 U346 ( .A1(n200), .A2(n193), .ZN(n359) );
  XOR2_X1 U347 ( .A(n263), .B(a[4]), .Z(n357) );
  INV_X1 U348 ( .A(n30), .ZN(n28) );
  INV_X1 U349 ( .A(n64), .ZN(n103) );
  INV_X1 U350 ( .A(n31), .ZN(n29) );
  INV_X1 U351 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U352 ( .A1(n52), .A2(n32), .ZN(n30) );
  INV_X1 U353 ( .A(n75), .ZN(n74) );
  NAND2_X1 U354 ( .A1(n356), .A2(n82), .ZN(n13) );
  XNOR2_X1 U355 ( .A(n16), .B(n306), .ZN(product[2]) );
  NAND2_X1 U356 ( .A1(n359), .A2(n94), .ZN(n16) );
  NAND2_X1 U357 ( .A1(n312), .A2(n62), .ZN(n8) );
  NAND2_X1 U358 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U359 ( .A(n34), .ZN(n99) );
  INV_X1 U360 ( .A(n82), .ZN(n80) );
  XNOR2_X1 U361 ( .A(n12), .B(n358), .ZN(product[6]) );
  INV_X1 U362 ( .A(n346), .ZN(n358) );
  XNOR2_X1 U363 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U364 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U365 ( .A(n23), .ZN(n98) );
  XNOR2_X1 U366 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U367 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U368 ( .A(n41), .ZN(n100) );
  NAND2_X1 U369 ( .A1(n329), .A2(n70), .ZN(n10) );
  OAI21_X1 U370 ( .B1(n76), .B2(n345), .A(n77), .ZN(n75) );
  AOI21_X1 U371 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U372 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U373 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U374 ( .A1(n52), .A2(n51), .ZN(n7) );
  XOR2_X1 U375 ( .A(n74), .B(n11), .Z(product[7]) );
  NAND2_X1 U376 ( .A1(n105), .A2(n73), .ZN(n11) );
  INV_X1 U377 ( .A(n72), .ZN(n105) );
  NOR2_X1 U378 ( .A1(n41), .A2(n34), .ZN(n32) );
  OAI21_X1 U379 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  OAI21_X1 U380 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  INV_X1 U381 ( .A(n50), .ZN(n52) );
  AOI21_X1 U382 ( .B1(n359), .B2(n306), .A(n92), .ZN(n90) );
  INV_X1 U383 ( .A(n94), .ZN(n92) );
  NAND2_X1 U384 ( .A1(n125), .A2(n130), .ZN(n65) );
  OAI21_X1 U385 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  NOR2_X1 U386 ( .A1(n30), .A2(n23), .ZN(n21) );
  INV_X1 U387 ( .A(n51), .ZN(n53) );
  NAND2_X1 U388 ( .A1(n131), .A2(n136), .ZN(n70) );
  NOR2_X1 U389 ( .A1(n50), .A2(n41), .ZN(n39) );
  XOR2_X1 U390 ( .A(n15), .B(n90), .Z(product[3]) );
  NOR2_X1 U391 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U392 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U393 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U394 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U395 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U396 ( .A(n84), .ZN(n108) );
  NOR2_X1 U397 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U398 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U399 ( .A(n112), .ZN(n113) );
  NAND2_X1 U400 ( .A1(n170), .A2(n112), .ZN(n24) );
  AND2_X1 U401 ( .A1(n363), .A2(n161), .ZN(n193) );
  NAND2_X1 U402 ( .A1(n116), .A2(n115), .ZN(n44) );
  NAND2_X1 U403 ( .A1(n200), .A2(n193), .ZN(n94) );
  NAND2_X1 U404 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U405 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U406 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U407 ( .A1(n147), .A2(n150), .ZN(n82) );
  NAND2_X1 U408 ( .A1(n143), .A2(n146), .ZN(n77) );
  INV_X1 U409 ( .A(n157), .ZN(n178) );
  OAI22_X1 U410 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  AND2_X1 U411 ( .A1(n363), .A2(n158), .ZN(n185) );
  OAI22_X1 U412 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  INV_X1 U413 ( .A(n118), .ZN(n119) );
  OR2_X1 U414 ( .A1(n363), .A2(n259), .ZN(n219) );
  AND2_X1 U415 ( .A1(n330), .A2(n97), .ZN(product[1]) );
  INV_X1 U416 ( .A(n163), .ZN(n194) );
  OAI22_X1 U417 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  OAI22_X1 U418 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  AND2_X1 U419 ( .A1(n363), .A2(n343), .ZN(n177) );
  OAI22_X1 U420 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  NOR2_X1 U421 ( .A1(n151), .A2(n152), .ZN(n84) );
  NOR2_X1 U422 ( .A1(n153), .A2(n168), .ZN(n88) );
  INV_X1 U423 ( .A(n154), .ZN(n170) );
  NAND2_X1 U424 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U425 ( .A1(n363), .A2(n258), .ZN(n210) );
  OR2_X1 U426 ( .A1(n363), .A2(n260), .ZN(n228) );
  OAI22_X1 U427 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U428 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  NAND2_X1 U429 ( .A1(n361), .A2(n333), .ZN(n252) );
  AND2_X1 U430 ( .A1(n363), .A2(n164), .ZN(product[0]) );
  XNOR2_X1 U431 ( .A(n264), .B(a[4]), .ZN(n255) );
  NAND2_X2 U432 ( .A1(n249), .A2(n273), .ZN(n253) );
  BUF_X1 U433 ( .A(n256), .Z(n361) );
  XNOR2_X1 U434 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U435 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U436 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U437 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U438 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U439 ( .A(n318), .B(n262), .ZN(n206) );
  XNOR2_X1 U440 ( .A(n262), .B(n363), .ZN(n209) );
  INV_X1 U441 ( .A(n262), .ZN(n258) );
  XNOR2_X1 U442 ( .A(b[1]), .B(n262), .ZN(n208) );
  NAND2_X1 U443 ( .A1(n308), .A2(n21), .ZN(n19) );
  NAND2_X1 U444 ( .A1(n308), .A2(n28), .ZN(n26) );
  XNOR2_X1 U445 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U446 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U447 ( .A1(n308), .A2(n39), .ZN(n37) );
  INV_X1 U448 ( .A(n3), .ZN(n57) );
  INV_X1 U449 ( .A(n88), .ZN(n109) );
  OAI21_X1 U450 ( .B1(n338), .B2(n73), .A(n70), .ZN(n68) );
  NOR2_X1 U451 ( .A1(n69), .A2(n72), .ZN(n67) );
  XOR2_X1 U452 ( .A(n14), .B(n314), .Z(product[4]) );
  AOI21_X1 U453 ( .B1(n337), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U454 ( .B1(n337), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U455 ( .A(n337), .ZN(n58) );
  AOI21_X1 U456 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U457 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  INV_X1 U458 ( .A(n128), .ZN(n129) );
  INV_X1 U459 ( .A(n87), .ZN(n86) );
  XNOR2_X1 U460 ( .A(n13), .B(n304), .ZN(product[5]) );
  NAND2_X1 U461 ( .A1(n109), .A2(n316), .ZN(n15) );
  OAI21_X1 U462 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  INV_X1 U463 ( .A(n160), .ZN(n186) );
  XNOR2_X1 U464 ( .A(n63), .B(n8), .ZN(product[10]) );
  XNOR2_X1 U465 ( .A(n71), .B(n10), .ZN(product[8]) );
  OAI21_X1 U466 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  OAI21_X1 U467 ( .B1(n354), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U468 ( .B1(n351), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U469 ( .B1(n351), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U470 ( .B1(n354), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U471 ( .B1(n351), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U472 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  XNOR2_X1 U473 ( .A(n264), .B(b[3]), .ZN(n224) );
  INV_X1 U474 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U475 ( .A(n264), .B(b[4]), .ZN(n223) );
  XNOR2_X1 U476 ( .A(b[5]), .B(n313), .ZN(n222) );
  XNOR2_X1 U477 ( .A(b[2]), .B(n332), .ZN(n225) );
  XNOR2_X1 U478 ( .A(b[6]), .B(n332), .ZN(n221) );
  XNOR2_X1 U479 ( .A(n303), .B(n363), .ZN(n227) );
  XNOR2_X1 U480 ( .A(b[7]), .B(n309), .ZN(n220) );
  XNOR2_X1 U481 ( .A(b[1]), .B(n303), .ZN(n226) );
  XOR2_X1 U482 ( .A(n264), .B(a[2]), .Z(n248) );
  OAI22_X1 U483 ( .A1(n341), .A2(n217), .B1(n216), .B2(n347), .ZN(n183) );
  OAI22_X1 U484 ( .A1(n342), .A2(n212), .B1(n211), .B2(n347), .ZN(n118) );
  OAI22_X1 U485 ( .A1(n211), .A2(n341), .B1(n211), .B2(n347), .ZN(n157) );
  OAI22_X1 U486 ( .A1(n342), .A2(n214), .B1(n213), .B2(n347), .ZN(n180) );
  OAI22_X1 U487 ( .A1(n341), .A2(n213), .B1(n212), .B2(n347), .ZN(n179) );
  OAI22_X1 U488 ( .A1(n341), .A2(n216), .B1(n215), .B2(n347), .ZN(n182) );
  OAI22_X1 U489 ( .A1(n342), .A2(n215), .B1(n214), .B2(n347), .ZN(n181) );
  INV_X1 U490 ( .A(n347), .ZN(n158) );
  OAI22_X1 U491 ( .A1(n323), .A2(n259), .B1(n219), .B2(n347), .ZN(n167) );
  OAI22_X1 U492 ( .A1(n323), .A2(n218), .B1(n217), .B2(n347), .ZN(n184) );
  OAI22_X1 U493 ( .A1(n353), .A2(n221), .B1(n220), .B2(n311), .ZN(n128) );
  OAI22_X1 U494 ( .A1(n305), .A2(n260), .B1(n228), .B2(n311), .ZN(n168) );
  OAI22_X1 U495 ( .A1(n353), .A2(n225), .B1(n315), .B2(n311), .ZN(n190) );
  OAI22_X1 U496 ( .A1(n252), .A2(n224), .B1(n223), .B2(n362), .ZN(n189) );
  OAI22_X1 U497 ( .A1(n305), .A2(n222), .B1(n221), .B2(n311), .ZN(n187) );
  OAI22_X1 U498 ( .A1(n220), .A2(n353), .B1(n220), .B2(n311), .ZN(n160) );
  OAI22_X1 U499 ( .A1(n353), .A2(n223), .B1(n222), .B2(n311), .ZN(n188) );
  OAI22_X1 U500 ( .A1(n353), .A2(n226), .B1(n225), .B2(n311), .ZN(n191) );
  XNOR2_X1 U501 ( .A(b[5]), .B(n335), .ZN(n231) );
  OAI22_X1 U502 ( .A1(n252), .A2(n227), .B1(n226), .B2(n362), .ZN(n192) );
  XNOR2_X1 U503 ( .A(b[6]), .B(n334), .ZN(n230) );
  INV_X1 U504 ( .A(n362), .ZN(n161) );
  XNOR2_X1 U505 ( .A(b[4]), .B(n335), .ZN(n232) );
  XNOR2_X1 U506 ( .A(n334), .B(b[3]), .ZN(n233) );
  XNOR2_X1 U507 ( .A(n335), .B(n363), .ZN(n236) );
  XNOR2_X1 U508 ( .A(b[2]), .B(n335), .ZN(n234) );
  XNOR2_X1 U509 ( .A(b[7]), .B(n334), .ZN(n229) );
  INV_X1 U510 ( .A(n334), .ZN(n261) );
  XNOR2_X1 U511 ( .A(b[1]), .B(n334), .ZN(n235) );
  XOR2_X1 U512 ( .A(n265), .B(n164), .Z(n249) );
  XNOR2_X1 U513 ( .A(n265), .B(a[2]), .ZN(n256) );
  OAI22_X1 U514 ( .A1(n202), .A2(n339), .B1(n202), .B2(n349), .ZN(n154) );
  OAI22_X1 U515 ( .A1(n339), .A2(n203), .B1(n202), .B2(n350), .ZN(n112) );
  OAI22_X1 U516 ( .A1(n339), .A2(n206), .B1(n205), .B2(n349), .ZN(n173) );
  OAI22_X1 U517 ( .A1(n339), .A2(n205), .B1(n204), .B2(n349), .ZN(n172) );
  OAI22_X1 U518 ( .A1(n339), .A2(n204), .B1(n203), .B2(n350), .ZN(n171) );
  OAI22_X1 U519 ( .A1(n339), .A2(n207), .B1(n206), .B2(n350), .ZN(n174) );
  XNOR2_X1 U520 ( .A(b[7]), .B(n340), .ZN(n211) );
  OAI22_X1 U521 ( .A1(n339), .A2(n208), .B1(n207), .B2(n349), .ZN(n175) );
  XNOR2_X1 U522 ( .A(b[6]), .B(n340), .ZN(n212) );
  XNOR2_X1 U523 ( .A(b[5]), .B(n340), .ZN(n213) );
  OAI22_X1 U524 ( .A1(n250), .A2(n258), .B1(n210), .B2(n350), .ZN(n166) );
  OAI22_X1 U525 ( .A1(n250), .A2(n209), .B1(n208), .B2(n349), .ZN(n176) );
  XNOR2_X1 U526 ( .A(b[2]), .B(n328), .ZN(n216) );
  XNOR2_X1 U527 ( .A(b[4]), .B(n327), .ZN(n214) );
  XNOR2_X1 U528 ( .A(n327), .B(n363), .ZN(n218) );
  INV_X1 U529 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U530 ( .A(b[1]), .B(n263), .ZN(n217) );
  NAND2_X1 U531 ( .A1(n153), .A2(n168), .ZN(n89) );
  INV_X2 U532 ( .A(n164), .ZN(n273) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n12, n13, n14, n15, n16, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50,
         n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102, n103,
         n104, n109, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n157, n158, n160, n161, n163, n164, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n245, n246, n249, n250, n251, n252, n253, n254,
         n255, n256, n258, n259, n260, n262, n263, n264, n265, n273, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n369, n370,
         n371, n372, n373;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n128), .B(n179), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  XNOR2_X2 U268 ( .A(n263), .B(a[6]), .ZN(n254) );
  CLKBUF_X3 U269 ( .A(n263), .Z(n351) );
  CLKBUF_X1 U270 ( .A(n319), .Z(n303) );
  BUF_X1 U271 ( .A(n75), .Z(n308) );
  OAI21_X1 U272 ( .B1(n84), .B2(n86), .A(n85), .ZN(n304) );
  AND2_X1 U273 ( .A1(n52), .A2(n102), .ZN(n305) );
  INV_X1 U274 ( .A(n58), .ZN(n306) );
  OR2_X1 U275 ( .A1(n137), .A2(n142), .ZN(n307) );
  BUF_X1 U276 ( .A(n75), .Z(n332) );
  CLKBUF_X1 U277 ( .A(n252), .Z(n309) );
  BUF_X1 U278 ( .A(n256), .Z(n371) );
  XNOR2_X1 U279 ( .A(n74), .B(n310), .ZN(product[7]) );
  AND2_X1 U280 ( .A1(n307), .A2(n73), .ZN(n310) );
  OR2_X1 U281 ( .A1(n151), .A2(n152), .ZN(n311) );
  XOR2_X1 U282 ( .A(n148), .B(n183), .Z(n312) );
  XOR2_X1 U283 ( .A(n145), .B(n312), .Z(n143) );
  NAND2_X1 U284 ( .A1(n145), .A2(n148), .ZN(n313) );
  NAND2_X1 U285 ( .A1(n145), .A2(n183), .ZN(n314) );
  NAND2_X1 U286 ( .A1(n148), .A2(n183), .ZN(n315) );
  NAND3_X1 U287 ( .A1(n313), .A2(n314), .A3(n315), .ZN(n142) );
  BUF_X1 U288 ( .A(n255), .Z(n372) );
  OAI21_X1 U289 ( .B1(n73), .B2(n69), .A(n70), .ZN(n316) );
  XNOR2_X1 U290 ( .A(n263), .B(a[6]), .ZN(n363) );
  INV_X1 U291 ( .A(n259), .ZN(n317) );
  NOR2_X2 U292 ( .A1(n131), .A2(n136), .ZN(n69) );
  BUF_X1 U293 ( .A(n264), .Z(n339) );
  CLKBUF_X3 U294 ( .A(n337), .Z(n318) );
  OR2_X2 U295 ( .A1(n147), .A2(n150), .ZN(n367) );
  BUF_X1 U296 ( .A(n265), .Z(n333) );
  BUF_X1 U297 ( .A(n256), .Z(n350) );
  NAND2_X1 U298 ( .A1(n364), .A2(n337), .ZN(n319) );
  NAND2_X1 U299 ( .A1(n364), .A2(n337), .ZN(n251) );
  XNOR2_X1 U300 ( .A(n133), .B(n320), .ZN(n131) );
  XNOR2_X1 U301 ( .A(n138), .B(n135), .ZN(n320) );
  CLKBUF_X1 U302 ( .A(n362), .Z(n321) );
  XNOR2_X1 U303 ( .A(n187), .B(n175), .ZN(n135) );
  NAND2_X1 U304 ( .A1(n355), .A2(n356), .ZN(n322) );
  CLKBUF_X1 U305 ( .A(n265), .Z(n323) );
  NAND2_X1 U306 ( .A1(n133), .A2(n138), .ZN(n324) );
  NAND2_X1 U307 ( .A1(n133), .A2(n135), .ZN(n325) );
  NAND2_X1 U308 ( .A1(n138), .A2(n135), .ZN(n326) );
  NAND3_X1 U309 ( .A1(n324), .A2(n325), .A3(n326), .ZN(n130) );
  NAND2_X1 U310 ( .A1(n262), .A2(n373), .ZN(n328) );
  NAND2_X1 U311 ( .A1(n258), .A2(n327), .ZN(n329) );
  NAND2_X1 U312 ( .A1(n328), .A2(n329), .ZN(n209) );
  INV_X1 U313 ( .A(n373), .ZN(n327) );
  NOR2_X1 U314 ( .A1(n137), .A2(n142), .ZN(n72) );
  NOR2_X1 U315 ( .A1(n121), .A2(n124), .ZN(n61) );
  OR2_X1 U316 ( .A1(n201), .A2(n169), .ZN(n330) );
  XNOR2_X1 U317 ( .A(n362), .B(n331), .ZN(product[9]) );
  AND2_X1 U318 ( .A1(n103), .A2(n65), .ZN(n331) );
  BUF_X1 U319 ( .A(n256), .Z(n334) );
  BUF_X2 U320 ( .A(n339), .Z(n335) );
  CLKBUF_X1 U321 ( .A(n263), .Z(n336) );
  XNOR2_X1 U322 ( .A(n339), .B(a[4]), .ZN(n337) );
  OR2_X1 U323 ( .A1(n143), .A2(n146), .ZN(n338) );
  INV_X1 U324 ( .A(n342), .ZN(n82) );
  AND2_X1 U325 ( .A1(n147), .A2(n150), .ZN(n342) );
  CLKBUF_X1 U326 ( .A(n264), .Z(n370) );
  NAND2_X1 U327 ( .A1(n246), .A2(n363), .ZN(n340) );
  NAND2_X1 U328 ( .A1(n246), .A2(n254), .ZN(n341) );
  NAND2_X1 U329 ( .A1(n246), .A2(n363), .ZN(n250) );
  NAND2_X1 U330 ( .A1(a[6]), .A2(n344), .ZN(n345) );
  NAND2_X1 U331 ( .A1(n343), .A2(n262), .ZN(n346) );
  NAND2_X1 U332 ( .A1(n345), .A2(n346), .ZN(n246) );
  INV_X1 U333 ( .A(a[6]), .ZN(n343) );
  INV_X1 U334 ( .A(n262), .ZN(n344) );
  AOI21_X2 U335 ( .B1(n67), .B2(n332), .A(n316), .ZN(n362) );
  CLKBUF_X1 U336 ( .A(n89), .Z(n347) );
  NAND2_X1 U337 ( .A1(n249), .A2(n273), .ZN(n348) );
  NAND2_X1 U338 ( .A1(n322), .A2(n273), .ZN(n349) );
  NAND2_X1 U339 ( .A1(n322), .A2(n273), .ZN(n253) );
  BUF_X1 U340 ( .A(b[3]), .Z(n352) );
  BUF_X1 U341 ( .A(n264), .Z(n369) );
  BUF_X2 U342 ( .A(n245), .Z(n373) );
  NAND2_X1 U343 ( .A1(n265), .A2(n354), .ZN(n355) );
  NAND2_X1 U344 ( .A1(n353), .A2(n164), .ZN(n356) );
  NAND2_X1 U345 ( .A1(n355), .A2(n356), .ZN(n249) );
  INV_X1 U346 ( .A(n265), .ZN(n353) );
  INV_X1 U347 ( .A(n164), .ZN(n354) );
  NAND2_X1 U348 ( .A1(n365), .A2(n334), .ZN(n357) );
  NAND2_X1 U349 ( .A1(n359), .A2(n334), .ZN(n358) );
  XOR2_X1 U350 ( .A(n370), .B(a[2]), .Z(n359) );
  NAND2_X1 U351 ( .A1(n365), .A2(n256), .ZN(n252) );
  CLKBUF_X1 U352 ( .A(n304), .Z(n360) );
  AOI21_X1 U353 ( .B1(n367), .B2(n304), .A(n342), .ZN(n361) );
  AOI21_X1 U354 ( .B1(n67), .B2(n308), .A(n68), .ZN(n1) );
  NOR2_X1 U355 ( .A1(n64), .A2(n61), .ZN(n3) );
  NOR2_X1 U356 ( .A1(n125), .A2(n130), .ZN(n64) );
  NAND2_X1 U357 ( .A1(n137), .A2(n142), .ZN(n73) );
  XOR2_X1 U358 ( .A(n263), .B(a[4]), .Z(n364) );
  XOR2_X1 U359 ( .A(n369), .B(a[2]), .Z(n365) );
  INV_X1 U360 ( .A(n30), .ZN(n28) );
  INV_X1 U361 ( .A(n64), .ZN(n103) );
  INV_X1 U362 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U363 ( .A1(n3), .A2(n21), .ZN(n19) );
  AOI21_X1 U364 ( .B1(n306), .B2(n21), .A(n22), .ZN(n20) );
  INV_X1 U365 ( .A(n31), .ZN(n29) );
  INV_X1 U366 ( .A(n75), .ZN(n74) );
  NAND2_X1 U367 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U368 ( .A1(n3), .A2(n39), .ZN(n37) );
  INV_X1 U369 ( .A(n2), .ZN(n58) );
  NAND2_X1 U370 ( .A1(n109), .A2(n347), .ZN(n15) );
  INV_X1 U371 ( .A(n88), .ZN(n109) );
  NAND2_X1 U372 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U373 ( .A(n23), .ZN(n98) );
  XNOR2_X1 U374 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U375 ( .A1(n366), .A2(n94), .ZN(n16) );
  NAND2_X1 U376 ( .A1(n52), .A2(n51), .ZN(n7) );
  INV_X1 U377 ( .A(n3), .ZN(n57) );
  NAND2_X1 U378 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U379 ( .A(n41), .ZN(n100) );
  OAI21_X1 U380 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  INV_X1 U381 ( .A(n94), .ZN(n92) );
  XNOR2_X1 U382 ( .A(n13), .B(n360), .ZN(product[5]) );
  NAND2_X1 U383 ( .A1(n367), .A2(n82), .ZN(n13) );
  NAND2_X1 U384 ( .A1(n338), .A2(n77), .ZN(n12) );
  XNOR2_X1 U385 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U386 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U387 ( .A(n61), .ZN(n102) );
  OAI21_X1 U388 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  AOI21_X1 U389 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U390 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U391 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U392 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U393 ( .A(n34), .ZN(n99) );
  NOR2_X1 U394 ( .A1(n30), .A2(n23), .ZN(n21) );
  XOR2_X1 U395 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U396 ( .A1(n311), .A2(n85), .ZN(n14) );
  NOR2_X1 U397 ( .A1(n50), .A2(n41), .ZN(n39) );
  NOR2_X1 U398 ( .A1(n41), .A2(n34), .ZN(n32) );
  INV_X1 U399 ( .A(n50), .ZN(n52) );
  XNOR2_X1 U400 ( .A(n71), .B(n10), .ZN(product[8]) );
  NAND2_X1 U401 ( .A1(n104), .A2(n70), .ZN(n10) );
  OAI21_X1 U402 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  INV_X1 U403 ( .A(n69), .ZN(n104) );
  OAI21_X1 U404 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  NAND2_X1 U405 ( .A1(n125), .A2(n130), .ZN(n65) );
  AOI21_X1 U406 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U407 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  INV_X1 U408 ( .A(n51), .ZN(n53) );
  NAND2_X1 U409 ( .A1(n131), .A2(n136), .ZN(n70) );
  INV_X1 U410 ( .A(n87), .ZN(n86) );
  NOR2_X1 U411 ( .A1(n116), .A2(n115), .ZN(n41) );
  OR2_X1 U412 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U413 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U414 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U415 ( .A(n112), .ZN(n113) );
  NOR2_X1 U416 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U417 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U418 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U419 ( .A1(n151), .A2(n152), .ZN(n84) );
  NAND2_X1 U420 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U421 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U422 ( .A1(n121), .A2(n124), .ZN(n62) );
  INV_X1 U423 ( .A(n97), .ZN(n95) );
  NAND2_X1 U424 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U425 ( .A1(n200), .A2(n193), .ZN(n366) );
  NAND2_X1 U426 ( .A1(n143), .A2(n146), .ZN(n77) );
  AND2_X1 U427 ( .A1(n373), .A2(n161), .ZN(n193) );
  OR2_X1 U428 ( .A1(n373), .A2(n260), .ZN(n228) );
  INV_X1 U429 ( .A(n157), .ZN(n178) );
  AND2_X1 U430 ( .A1(n373), .A2(n158), .ZN(n185) );
  OAI22_X1 U431 ( .A1(n349), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  INV_X1 U432 ( .A(n118), .ZN(n119) );
  OAI22_X1 U433 ( .A1(n234), .A2(n348), .B1(n233), .B2(n273), .ZN(n199) );
  OR2_X1 U434 ( .A1(n373), .A2(n259), .ZN(n219) );
  OAI22_X1 U435 ( .A1(n349), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  AND2_X1 U436 ( .A1(n330), .A2(n97), .ZN(product[1]) );
  INV_X1 U437 ( .A(n163), .ZN(n194) );
  OAI22_X1 U438 ( .A1(n229), .A2(n349), .B1(n229), .B2(n273), .ZN(n163) );
  INV_X1 U439 ( .A(n128), .ZN(n129) );
  AND2_X1 U440 ( .A1(n373), .A2(n155), .ZN(n177) );
  OAI22_X1 U441 ( .A1(n348), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U442 ( .A1(n349), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  INV_X1 U443 ( .A(n154), .ZN(n170) );
  OR2_X1 U444 ( .A1(n373), .A2(n258), .ZN(n210) );
  INV_X1 U445 ( .A(n160), .ZN(n186) );
  OAI22_X1 U446 ( .A1(n253), .A2(n353), .B1(n237), .B2(n273), .ZN(n169) );
  OR2_X1 U447 ( .A1(n373), .A2(n353), .ZN(n237) );
  XNOR2_X1 U448 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U449 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U450 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U451 ( .A(b[6]), .B(n262), .ZN(n203) );
  INV_X1 U452 ( .A(n262), .ZN(n258) );
  AND2_X1 U453 ( .A1(n245), .A2(n164), .ZN(product[0]) );
  XOR2_X1 U454 ( .A(n15), .B(n90), .Z(product[3]) );
  NOR2_X1 U455 ( .A1(n143), .A2(n146), .ZN(n76) );
  XNOR2_X1 U456 ( .A(n265), .B(a[2]), .ZN(n256) );
  XNOR2_X1 U457 ( .A(n369), .B(a[4]), .ZN(n255) );
  XNOR2_X1 U458 ( .A(n56), .B(n7), .ZN(product[11]) );
  INV_X1 U459 ( .A(n335), .ZN(n260) );
  XNOR2_X1 U460 ( .A(n370), .B(b[5]), .ZN(n222) );
  XNOR2_X1 U461 ( .A(n335), .B(n373), .ZN(n227) );
  XNOR2_X1 U462 ( .A(b[4]), .B(n335), .ZN(n223) );
  XNOR2_X1 U463 ( .A(n370), .B(b[6]), .ZN(n221) );
  NOR2_X1 U464 ( .A1(n153), .A2(n168), .ZN(n88) );
  XNOR2_X1 U465 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U466 ( .A1(n305), .A2(n103), .ZN(n46) );
  AOI21_X1 U467 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  OAI22_X1 U468 ( .A1(n202), .A2(n340), .B1(n202), .B2(n254), .ZN(n154) );
  OAI22_X1 U469 ( .A1(n341), .A2(n203), .B1(n254), .B2(n202), .ZN(n112) );
  OAI22_X1 U470 ( .A1(n340), .A2(n205), .B1(n254), .B2(n204), .ZN(n172) );
  OAI22_X1 U471 ( .A1(n340), .A2(n206), .B1(n254), .B2(n205), .ZN(n173) );
  OAI22_X1 U472 ( .A1(n341), .A2(n204), .B1(n254), .B2(n203), .ZN(n171) );
  OAI22_X1 U473 ( .A1(n341), .A2(n208), .B1(n254), .B2(n207), .ZN(n175) );
  XNOR2_X1 U474 ( .A(n351), .B(b[7]), .ZN(n211) );
  OAI22_X1 U475 ( .A1(n340), .A2(n207), .B1(n254), .B2(n206), .ZN(n174) );
  INV_X1 U476 ( .A(n363), .ZN(n155) );
  OAI22_X1 U477 ( .A1(n250), .A2(n209), .B1(n254), .B2(n208), .ZN(n176) );
  OAI22_X1 U478 ( .A1(n250), .A2(n258), .B1(n210), .B2(n363), .ZN(n166) );
  XNOR2_X1 U479 ( .A(n317), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U480 ( .A(n351), .B(n373), .ZN(n218) );
  XNOR2_X1 U481 ( .A(n351), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U482 ( .A(n351), .B(b[6]), .ZN(n212) );
  INV_X1 U483 ( .A(n263), .ZN(n259) );
  NAND2_X1 U484 ( .A1(n200), .A2(n193), .ZN(n94) );
  AOI21_X1 U485 ( .B1(n366), .B2(n95), .A(n92), .ZN(n90) );
  OAI21_X1 U486 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  OAI22_X1 U487 ( .A1(n349), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  XNOR2_X1 U488 ( .A(n25), .B(n4), .ZN(product[14]) );
  AOI21_X1 U489 ( .B1(n306), .B2(n28), .A(n29), .ZN(n27) );
  XNOR2_X1 U490 ( .A(n370), .B(b[7]), .ZN(n220) );
  OAI21_X1 U491 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  XNOR2_X1 U492 ( .A(n351), .B(n352), .ZN(n215) );
  XNOR2_X1 U493 ( .A(n335), .B(b[3]), .ZN(n224) );
  XNOR2_X1 U494 ( .A(n352), .B(n262), .ZN(n206) );
  XNOR2_X1 U495 ( .A(n336), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U496 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U497 ( .A(n335), .B(b[2]), .ZN(n225) );
  XNOR2_X1 U498 ( .A(b[1]), .B(n262), .ZN(n208) );
  XNOR2_X1 U499 ( .A(n336), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U500 ( .A(n370), .B(b[1]), .ZN(n226) );
  OAI21_X1 U501 ( .B1(n73), .B2(n69), .A(n70), .ZN(n68) );
  NOR2_X1 U502 ( .A1(n69), .A2(n72), .ZN(n67) );
  NAND2_X1 U503 ( .A1(n3), .A2(n28), .ZN(n26) );
  NAND2_X1 U504 ( .A1(n201), .A2(n169), .ZN(n97) );
  AOI21_X1 U505 ( .B1(n367), .B2(n83), .A(n342), .ZN(n78) );
  XOR2_X1 U506 ( .A(n12), .B(n361), .Z(product[6]) );
  OAI22_X1 U507 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  NAND2_X1 U508 ( .A1(n153), .A2(n168), .ZN(n89) );
  OAI22_X1 U509 ( .A1(n319), .A2(n217), .B1(n216), .B2(n318), .ZN(n183) );
  OAI22_X1 U510 ( .A1(n319), .A2(n216), .B1(n215), .B2(n318), .ZN(n182) );
  OAI22_X1 U511 ( .A1(n303), .A2(n212), .B1(n211), .B2(n318), .ZN(n118) );
  OAI22_X1 U512 ( .A1(n319), .A2(n215), .B1(n214), .B2(n318), .ZN(n181) );
  OAI22_X1 U513 ( .A1(n319), .A2(n214), .B1(n213), .B2(n318), .ZN(n180) );
  OAI22_X1 U514 ( .A1(n211), .A2(n303), .B1(n211), .B2(n318), .ZN(n157) );
  OAI22_X1 U515 ( .A1(n319), .A2(n213), .B1(n212), .B2(n318), .ZN(n179) );
  INV_X1 U516 ( .A(n372), .ZN(n158) );
  OAI22_X1 U517 ( .A1(n251), .A2(n259), .B1(n219), .B2(n372), .ZN(n167) );
  OAI22_X1 U518 ( .A1(n251), .A2(n218), .B1(n217), .B2(n372), .ZN(n184) );
  OAI21_X1 U519 ( .B1(n321), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U520 ( .B1(n362), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U521 ( .B1(n321), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U522 ( .B1(n362), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U523 ( .B1(n362), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U524 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  OAI22_X1 U525 ( .A1(n357), .A2(n222), .B1(n221), .B2(n350), .ZN(n187) );
  OAI22_X1 U526 ( .A1(n309), .A2(n224), .B1(n223), .B2(n371), .ZN(n189) );
  OAI22_X1 U527 ( .A1(n357), .A2(n221), .B1(n220), .B2(n350), .ZN(n128) );
  OAI22_X1 U528 ( .A1(n358), .A2(n225), .B1(n224), .B2(n350), .ZN(n190) );
  OAI22_X1 U529 ( .A1(n358), .A2(n223), .B1(n222), .B2(n350), .ZN(n188) );
  OAI22_X1 U530 ( .A1(n220), .A2(n357), .B1(n220), .B2(n350), .ZN(n160) );
  OAI22_X1 U531 ( .A1(n358), .A2(n260), .B1(n228), .B2(n371), .ZN(n168) );
  OAI22_X1 U532 ( .A1(n358), .A2(n226), .B1(n225), .B2(n371), .ZN(n191) );
  XNOR2_X1 U533 ( .A(n323), .B(b[5]), .ZN(n231) );
  XNOR2_X1 U534 ( .A(n323), .B(b[6]), .ZN(n230) );
  OAI22_X1 U535 ( .A1(n252), .A2(n227), .B1(n226), .B2(n371), .ZN(n192) );
  INV_X1 U536 ( .A(n350), .ZN(n161) );
  XNOR2_X1 U537 ( .A(n333), .B(b[4]), .ZN(n232) );
  XNOR2_X1 U538 ( .A(n333), .B(b[7]), .ZN(n229) );
  XNOR2_X1 U539 ( .A(n333), .B(n373), .ZN(n236) );
  XNOR2_X1 U540 ( .A(n333), .B(b[3]), .ZN(n233) );
  XNOR2_X1 U541 ( .A(n333), .B(b[2]), .ZN(n234) );
  XNOR2_X1 U542 ( .A(n323), .B(b[1]), .ZN(n235) );
  INV_X2 U543 ( .A(n164), .ZN(n273) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_0_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n20, n21, n22, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n51, n52,
         n54, n56, n57, n58, n60, n62, n63, n64, n65, n66, n68, n70, n71, n72,
         n73, n74, n76, n78, n79, n80, n81, n82, n84, n86, n87, n89, n92, n93,
         n94, n95, n99, n101, n103, n160, n161, n162, n163, n164, n165, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183;

  AND2_X1 U125 ( .A1(A[14]), .A2(B[14]), .ZN(n160) );
  INV_X4 U126 ( .A(n160), .ZN(n26) );
  CLKBUF_X1 U127 ( .A(A[12]), .Z(n161) );
  BUF_X1 U128 ( .A(n169), .Z(n162) );
  CLKBUF_X1 U129 ( .A(n174), .Z(n163) );
  NOR2_X1 U130 ( .A1(B[10]), .A2(A[10]), .ZN(n42) );
  CLKBUF_X1 U131 ( .A(n170), .Z(n164) );
  BUF_X1 U132 ( .A(n33), .Z(n165) );
  INV_X1 U133 ( .A(n164), .ZN(n51) );
  AND2_X1 U134 ( .A1(n167), .A2(n89), .ZN(SUM[0]) );
  OR2_X1 U135 ( .A1(B[0]), .A2(A[0]), .ZN(n167) );
  XNOR2_X1 U136 ( .A(n44), .B(n168), .ZN(SUM[10]) );
  AND2_X1 U137 ( .A1(n95), .A2(n43), .ZN(n168) );
  OR2_X1 U138 ( .A1(B[9]), .A2(A[9]), .ZN(n169) );
  OR2_X1 U139 ( .A1(B[9]), .A2(A[9]), .ZN(n176) );
  AND2_X1 U140 ( .A1(B[9]), .A2(A[9]), .ZN(n170) );
  OR2_X2 U141 ( .A1(A[14]), .A2(B[14]), .ZN(n179) );
  AOI21_X1 U142 ( .B1(n45), .B2(n37), .A(n38), .ZN(n171) );
  AOI21_X1 U143 ( .B1(n45), .B2(n37), .A(n38), .ZN(n1) );
  NAND2_X1 U144 ( .A1(B[12]), .A2(n161), .ZN(n172) );
  INV_X1 U145 ( .A(n93), .ZN(n173) );
  NOR2_X1 U146 ( .A1(B[11]), .A2(A[11]), .ZN(n174) );
  NOR2_X1 U147 ( .A1(B[11]), .A2(A[11]), .ZN(n39) );
  NOR2_X1 U148 ( .A1(A[13]), .A2(B[13]), .ZN(n175) );
  INV_X1 U149 ( .A(n58), .ZN(n57) );
  INV_X1 U150 ( .A(n30), .ZN(n28) );
  OAI21_X1 U151 ( .B1(n64), .B2(n66), .A(n65), .ZN(n63) );
  AOI21_X1 U152 ( .B1(n71), .B2(n180), .A(n68), .ZN(n66) );
  NAND2_X1 U153 ( .A1(n93), .A2(n172), .ZN(n5) );
  INV_X1 U154 ( .A(n35), .ZN(n93) );
  NAND2_X1 U155 ( .A1(n92), .A2(n165), .ZN(n4) );
  NAND2_X1 U156 ( .A1(n179), .A2(n26), .ZN(n3) );
  AOI21_X1 U157 ( .B1(n178), .B2(n63), .A(n60), .ZN(n58) );
  INV_X1 U158 ( .A(n62), .ZN(n60) );
  NAND2_X1 U159 ( .A1(n99), .A2(n65), .ZN(n11) );
  INV_X1 U160 ( .A(n64), .ZN(n99) );
  XOR2_X1 U161 ( .A(n8), .B(n52), .Z(SUM[9]) );
  AOI21_X1 U162 ( .B1(n177), .B2(n57), .A(n54), .ZN(n52) );
  XNOR2_X1 U163 ( .A(n41), .B(n6), .ZN(SUM[11]) );
  NAND2_X1 U164 ( .A1(n94), .A2(n40), .ZN(n6) );
  INV_X1 U165 ( .A(n56), .ZN(n54) );
  XNOR2_X1 U166 ( .A(n9), .B(n57), .ZN(SUM[8]) );
  NAND2_X1 U167 ( .A1(n177), .A2(n56), .ZN(n9) );
  INV_X1 U168 ( .A(n42), .ZN(n95) );
  XNOR2_X1 U169 ( .A(n10), .B(n63), .ZN(SUM[7]) );
  NAND2_X1 U170 ( .A1(n178), .A2(n62), .ZN(n10) );
  NAND2_X1 U171 ( .A1(n180), .A2(n70), .ZN(n12) );
  NOR2_X1 U172 ( .A1(A[12]), .A2(B[12]), .ZN(n35) );
  OAI21_X1 U173 ( .B1(n72), .B2(n74), .A(n73), .ZN(n71) );
  OR2_X1 U174 ( .A1(B[8]), .A2(A[8]), .ZN(n177) );
  OR2_X1 U175 ( .A1(B[7]), .A2(A[7]), .ZN(n178) );
  AOI21_X1 U176 ( .B1(n182), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U177 ( .A(n78), .ZN(n76) );
  NAND2_X1 U178 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  NAND2_X1 U179 ( .A1(B[10]), .A2(A[10]), .ZN(n43) );
  NOR2_X1 U180 ( .A1(B[6]), .A2(A[6]), .ZN(n64) );
  NAND2_X1 U181 ( .A1(B[6]), .A2(A[6]), .ZN(n65) );
  OR2_X1 U182 ( .A1(B[5]), .A2(A[5]), .ZN(n180) );
  NAND2_X1 U183 ( .A1(n101), .A2(n73), .ZN(n13) );
  INV_X1 U184 ( .A(n72), .ZN(n101) );
  NAND2_X1 U185 ( .A1(n182), .A2(n78), .ZN(n14) );
  OR2_X1 U186 ( .A1(B[15]), .A2(A[15]), .ZN(n181) );
  OAI21_X1 U187 ( .B1(n82), .B2(n80), .A(n81), .ZN(n79) );
  OR2_X1 U188 ( .A1(B[3]), .A2(A[3]), .ZN(n182) );
  NAND2_X1 U189 ( .A1(B[4]), .A2(A[4]), .ZN(n73) );
  NOR2_X1 U190 ( .A1(B[4]), .A2(A[4]), .ZN(n72) );
  XOR2_X1 U191 ( .A(n15), .B(n82), .Z(SUM[2]) );
  NAND2_X1 U192 ( .A1(n103), .A2(n81), .ZN(n15) );
  INV_X1 U193 ( .A(n80), .ZN(n103) );
  INV_X1 U194 ( .A(n86), .ZN(n84) );
  XNOR2_X1 U195 ( .A(n16), .B(n87), .ZN(SUM[1]) );
  NAND2_X1 U196 ( .A1(n183), .A2(n86), .ZN(n16) );
  NAND2_X1 U197 ( .A1(B[2]), .A2(A[2]), .ZN(n81) );
  NAND2_X1 U198 ( .A1(B[1]), .A2(A[1]), .ZN(n86) );
  OR2_X1 U199 ( .A1(B[1]), .A2(A[1]), .ZN(n183) );
  INV_X1 U200 ( .A(n89), .ZN(n87) );
  NAND2_X1 U201 ( .A1(B[0]), .A2(A[0]), .ZN(n89) );
  XNOR2_X1 U202 ( .A(n14), .B(n79), .ZN(SUM[3]) );
  INV_X1 U203 ( .A(n70), .ZN(n68) );
  AOI21_X1 U204 ( .B1(n183), .B2(n87), .A(n84), .ZN(n82) );
  NOR2_X1 U205 ( .A1(B[2]), .A2(A[2]), .ZN(n80) );
  NAND2_X1 U206 ( .A1(B[5]), .A2(A[5]), .ZN(n70) );
  NAND2_X1 U207 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  NAND2_X1 U208 ( .A1(B[8]), .A2(A[8]), .ZN(n56) );
  XNOR2_X1 U209 ( .A(n12), .B(n71), .ZN(SUM[5]) );
  NAND2_X1 U210 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NOR2_X1 U211 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND2_X1 U212 ( .A1(n181), .A2(n19), .ZN(n2) );
  INV_X1 U213 ( .A(n31), .ZN(n29) );
  XOR2_X1 U214 ( .A(n13), .B(n74), .Z(SUM[4]) );
  XOR2_X1 U215 ( .A(n11), .B(n66), .Z(SUM[6]) );
  NAND2_X1 U216 ( .A1(B[3]), .A2(A[3]), .ZN(n78) );
  OAI21_X1 U217 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  INV_X1 U218 ( .A(n163), .ZN(n94) );
  NOR2_X1 U219 ( .A1(n174), .A2(n42), .ZN(n37) );
  OAI21_X1 U220 ( .B1(n39), .B2(n43), .A(n40), .ZN(n38) );
  NAND2_X1 U221 ( .A1(B[11]), .A2(A[11]), .ZN(n40) );
  INV_X1 U222 ( .A(n175), .ZN(n92) );
  NOR2_X1 U223 ( .A1(n175), .A2(n35), .ZN(n30) );
  OAI21_X1 U224 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U225 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  INV_X1 U226 ( .A(n45), .ZN(n44) );
  OAI21_X1 U227 ( .B1(n46), .B2(n58), .A(n47), .ZN(n45) );
  AOI21_X1 U228 ( .B1(n176), .B2(n54), .A(n170), .ZN(n47) );
  XNOR2_X1 U229 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U230 ( .A1(n30), .A2(n179), .ZN(n21) );
  AOI21_X1 U231 ( .B1(n31), .B2(n179), .A(n160), .ZN(n22) );
  XNOR2_X1 U232 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  NAND2_X1 U233 ( .A1(n162), .A2(n51), .ZN(n8) );
  NAND2_X1 U234 ( .A1(n169), .A2(n177), .ZN(n46) );
  XNOR2_X1 U235 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XOR2_X1 U236 ( .A(n171), .B(n5), .Z(SUM[12]) );
  OAI21_X1 U237 ( .B1(n21), .B2(n1), .A(n22), .ZN(n20) );
  OAI21_X1 U238 ( .B1(n171), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U239 ( .B1(n1), .B2(n173), .A(n172), .ZN(n34) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_0 ( .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;


  recursive_add_layer_INPUT_SCALE2_WIDTH16_0_DW01_add_2 add_56 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM(out) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_0_DW01_add_4 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n10, n11, n12, n13, n14, n15, n16, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n59, n60, n62, n64, n65, n66, n68, n70, n71, n72, n73,
         n74, n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89, n91, n93,
         n94, n95, n96, n98, n102, n104, n106, n162, n163, n164, n165, n166,
         n167, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184;

  CLKBUF_X1 U127 ( .A(n94), .Z(n162) );
  NOR2_X2 U128 ( .A1(B[11]), .A2(A[11]), .ZN(n42) );
  CLKBUF_X1 U129 ( .A(B[10]), .Z(n163) );
  CLKBUF_X1 U130 ( .A(n182), .Z(n164) );
  BUF_X1 U131 ( .A(n43), .Z(n165) );
  INV_X1 U132 ( .A(n166), .ZN(n59) );
  OR2_X2 U133 ( .A1(B[8]), .A2(A[8]), .ZN(n182) );
  AND2_X1 U134 ( .A1(B[8]), .A2(A[8]), .ZN(n166) );
  XNOR2_X1 U135 ( .A(n49), .B(n167), .ZN(SUM[10]) );
  NAND2_X1 U136 ( .A1(n175), .A2(n48), .ZN(n167) );
  AND2_X1 U137 ( .A1(n177), .A2(n91), .ZN(SUM[0]) );
  OR2_X1 U138 ( .A1(B[6]), .A2(A[6]), .ZN(n169) );
  XNOR2_X1 U139 ( .A(n1), .B(n170), .ZN(SUM[11]) );
  AND2_X1 U140 ( .A1(n96), .A2(n165), .ZN(n170) );
  INV_X1 U141 ( .A(n36), .ZN(n171) );
  OR2_X1 U142 ( .A1(n42), .A2(n173), .ZN(n172) );
  NOR2_X1 U143 ( .A1(A[12]), .A2(B[12]), .ZN(n173) );
  NOR2_X1 U144 ( .A1(B[9]), .A2(A[9]), .ZN(n50) );
  NOR2_X1 U145 ( .A1(A[10]), .A2(B[10]), .ZN(n174) );
  OR2_X1 U146 ( .A1(n163), .A2(A[10]), .ZN(n175) );
  CLKBUF_X1 U147 ( .A(n1), .Z(n176) );
  OR2_X1 U148 ( .A1(B[0]), .A2(A[0]), .ZN(n177) );
  XNOR2_X1 U149 ( .A(n52), .B(n178), .ZN(SUM[9]) );
  AND2_X1 U150 ( .A1(n98), .A2(n51), .ZN(n178) );
  INV_X1 U151 ( .A(n42), .ZN(n96) );
  NAND2_X1 U152 ( .A1(n102), .A2(n73), .ZN(n12) );
  INV_X1 U153 ( .A(n72), .ZN(n102) );
  NAND2_X1 U154 ( .A1(n93), .A2(n26), .ZN(n3) );
  INV_X1 U155 ( .A(n25), .ZN(n93) );
  XNOR2_X1 U156 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U157 ( .A1(n95), .A2(n40), .ZN(n5) );
  XNOR2_X1 U158 ( .A(n60), .B(n179), .ZN(SUM[8]) );
  AND2_X1 U159 ( .A1(n164), .A2(n59), .ZN(n179) );
  AOI21_X1 U160 ( .B1(n169), .B2(n71), .A(n68), .ZN(n66) );
  INV_X1 U161 ( .A(n70), .ZN(n68) );
  INV_X1 U162 ( .A(n33), .ZN(n31) );
  NAND2_X1 U163 ( .A1(n180), .A2(n19), .ZN(n2) );
  NAND2_X1 U164 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NAND2_X1 U165 ( .A1(n162), .A2(n33), .ZN(n4) );
  NOR2_X1 U166 ( .A1(n42), .A2(n39), .ZN(n37) );
  XNOR2_X1 U167 ( .A(n10), .B(n65), .ZN(SUM[7]) );
  NOR2_X1 U168 ( .A1(n32), .A2(n25), .ZN(n23) );
  INV_X1 U169 ( .A(n32), .ZN(n94) );
  OR2_X1 U170 ( .A1(B[15]), .A2(A[15]), .ZN(n180) );
  XNOR2_X1 U171 ( .A(n11), .B(n71), .ZN(SUM[6]) );
  NAND2_X1 U172 ( .A1(n169), .A2(n70), .ZN(n11) );
  NAND2_X1 U173 ( .A1(n184), .A2(n78), .ZN(n13) );
  INV_X1 U174 ( .A(n78), .ZN(n76) );
  INV_X1 U175 ( .A(n80), .ZN(n104) );
  NOR2_X1 U176 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  NOR2_X1 U177 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NOR2_X1 U178 ( .A1(B[10]), .A2(A[10]), .ZN(n47) );
  NOR2_X1 U179 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  OR2_X1 U180 ( .A1(B[2]), .A2(A[2]), .ZN(n181) );
  NAND2_X1 U181 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  NAND2_X1 U182 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U183 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  OR2_X1 U184 ( .A1(B[7]), .A2(A[7]), .ZN(n183) );
  OR2_X1 U185 ( .A1(B[4]), .A2(A[4]), .ZN(n184) );
  AOI21_X1 U186 ( .B1(n87), .B2(n181), .A(n84), .ZN(n82) );
  INV_X1 U187 ( .A(n86), .ZN(n84) );
  NAND2_X1 U188 ( .A1(B[3]), .A2(A[3]), .ZN(n81) );
  NOR2_X1 U189 ( .A1(B[3]), .A2(A[3]), .ZN(n80) );
  XNOR2_X1 U190 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U191 ( .A1(n181), .A2(n86), .ZN(n15) );
  XOR2_X1 U192 ( .A(n16), .B(n91), .Z(SUM[1]) );
  OAI21_X1 U193 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U194 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U195 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  NAND2_X1 U196 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  NAND2_X1 U197 ( .A1(A[9]), .A2(B[9]), .ZN(n51) );
  AOI21_X1 U198 ( .B1(n38), .B2(n94), .A(n31), .ZN(n29) );
  AOI21_X1 U199 ( .B1(n23), .B2(n171), .A(n24), .ZN(n22) );
  INV_X1 U200 ( .A(n38), .ZN(n36) );
  OAI21_X1 U201 ( .B1(n173), .B2(n43), .A(n40), .ZN(n38) );
  OAI21_X1 U202 ( .B1(n54), .B2(n66), .A(n55), .ZN(n53) );
  OAI21_X1 U203 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  AOI21_X1 U204 ( .B1(n184), .B2(n79), .A(n76), .ZN(n74) );
  XNOR2_X1 U205 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  NAND2_X1 U206 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  XOR2_X1 U207 ( .A(n14), .B(n82), .Z(SUM[3]) );
  NAND2_X1 U208 ( .A1(n104), .A2(n81), .ZN(n14) );
  NAND2_X1 U209 ( .A1(n37), .A2(n23), .ZN(n21) );
  NAND2_X1 U210 ( .A1(n37), .A2(n94), .ZN(n28) );
  NAND2_X1 U211 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  XOR2_X1 U212 ( .A(n12), .B(n74), .Z(SUM[5]) );
  NAND2_X1 U213 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  NAND2_X1 U214 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  NAND2_X1 U215 ( .A1(n106), .A2(n89), .ZN(n16) );
  INV_X1 U216 ( .A(n88), .ZN(n106) );
  INV_X1 U217 ( .A(n39), .ZN(n95) );
  OAI21_X1 U218 ( .B1(n47), .B2(n51), .A(n48), .ZN(n46) );
  INV_X1 U219 ( .A(n66), .ZN(n65) );
  NAND2_X1 U220 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  AOI21_X1 U221 ( .B1(n65), .B2(n183), .A(n62), .ZN(n60) );
  NAND2_X1 U222 ( .A1(n183), .A2(n64), .ZN(n10) );
  NAND2_X1 U223 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  AOI21_X1 U224 ( .B1(n182), .B2(n62), .A(n166), .ZN(n55) );
  INV_X1 U225 ( .A(n64), .ZN(n62) );
  OAI21_X1 U226 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  NOR2_X1 U227 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  OAI21_X1 U228 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  NAND2_X1 U229 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  XNOR2_X1 U230 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  XNOR2_X1 U231 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  INV_X1 U232 ( .A(n50), .ZN(n98) );
  NOR2_X1 U233 ( .A1(n174), .A2(n50), .ZN(n45) );
  XNOR2_X1 U234 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  OAI21_X1 U235 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  AOI21_X2 U236 ( .B1(n53), .B2(n45), .A(n46), .ZN(n1) );
  INV_X1 U237 ( .A(n53), .ZN(n52) );
  OAI21_X1 U238 ( .B1(n176), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U239 ( .B1(n28), .B2(n1), .A(n29), .ZN(n27) );
  OAI21_X1 U240 ( .B1(n1), .B2(n42), .A(n165), .ZN(n41) );
  OAI21_X1 U241 ( .B1(n1), .B2(n172), .A(n36), .ZN(n34) );
  NAND2_X1 U242 ( .A1(n182), .A2(n183), .ZN(n54) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_0_DW01_add_5 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n10, n11, n12, n13, n14, n15, n16, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51,
         n52, n53, n54, n55, n59, n60, n62, n64, n65, n66, n68, n70, n71, n72,
         n73, n74, n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89, n91,
         n93, n94, n96, n97, n102, n104, n106, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190;

  CLKBUF_X1 U127 ( .A(n183), .Z(n162) );
  NOR2_X1 U128 ( .A1(A[12]), .A2(B[12]), .ZN(n163) );
  CLKBUF_X1 U129 ( .A(A[12]), .Z(n164) );
  INV_X1 U130 ( .A(n96), .ZN(n165) );
  BUF_X1 U131 ( .A(n181), .Z(n166) );
  CLKBUF_X1 U132 ( .A(n38), .Z(n167) );
  OR2_X1 U133 ( .A1(B[8]), .A2(A[8]), .ZN(n168) );
  OR2_X1 U134 ( .A1(B[8]), .A2(A[8]), .ZN(n190) );
  OAI21_X1 U135 ( .B1(n51), .B2(n47), .A(n48), .ZN(n169) );
  INV_X1 U136 ( .A(n35), .ZN(n170) );
  AOI21_X1 U137 ( .B1(n182), .B2(n45), .A(n46), .ZN(n171) );
  AND2_X1 U138 ( .A1(n184), .A2(n91), .ZN(SUM[0]) );
  OR2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(n173) );
  OR2_X1 U140 ( .A1(B[9]), .A2(A[9]), .ZN(n174) );
  XNOR2_X1 U141 ( .A(n183), .B(n175), .ZN(SUM[11]) );
  AND2_X1 U142 ( .A1(n96), .A2(n43), .ZN(n175) );
  INV_X1 U143 ( .A(n176), .ZN(n59) );
  AND2_X1 U144 ( .A1(B[8]), .A2(A[8]), .ZN(n176) );
  CLKBUF_X1 U145 ( .A(n51), .Z(n177) );
  NOR2_X1 U146 ( .A1(A[9]), .A2(B[9]), .ZN(n178) );
  OR2_X1 U147 ( .A1(n164), .A2(B[12]), .ZN(n179) );
  XNOR2_X1 U148 ( .A(n180), .B(n52), .ZN(SUM[9]) );
  AND2_X1 U149 ( .A1(n174), .A2(n51), .ZN(n180) );
  NOR2_X1 U150 ( .A1(B[10]), .A2(A[10]), .ZN(n181) );
  NOR2_X1 U151 ( .A1(A[10]), .A2(B[10]), .ZN(n47) );
  BUF_X1 U152 ( .A(n53), .Z(n182) );
  AOI21_X1 U153 ( .B1(n182), .B2(n45), .A(n46), .ZN(n183) );
  AOI21_X1 U154 ( .B1(n182), .B2(n45), .A(n169), .ZN(n1) );
  NOR2_X1 U155 ( .A1(A[11]), .A2(B[11]), .ZN(n42) );
  OR2_X1 U156 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  INV_X1 U157 ( .A(n66), .ZN(n65) );
  XNOR2_X1 U158 ( .A(n11), .B(n71), .ZN(SUM[6]) );
  NAND2_X1 U159 ( .A1(n188), .A2(n70), .ZN(n11) );
  INV_X1 U160 ( .A(n42), .ZN(n96) );
  OAI21_X1 U161 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  XNOR2_X1 U162 ( .A(n49), .B(n7), .ZN(SUM[10]) );
  NAND2_X1 U163 ( .A1(n97), .A2(n48), .ZN(n7) );
  INV_X1 U164 ( .A(n166), .ZN(n97) );
  AOI21_X1 U165 ( .B1(n188), .B2(n71), .A(n68), .ZN(n66) );
  INV_X1 U166 ( .A(n70), .ZN(n68) );
  XNOR2_X1 U167 ( .A(n60), .B(n185), .ZN(SUM[8]) );
  AND2_X1 U168 ( .A1(n168), .A2(n59), .ZN(n185) );
  OAI21_X1 U169 ( .B1(n39), .B2(n43), .A(n40), .ZN(n38) );
  XOR2_X1 U170 ( .A(n12), .B(n74), .Z(SUM[5]) );
  INV_X1 U171 ( .A(n72), .ZN(n102) );
  INV_X1 U172 ( .A(n33), .ZN(n31) );
  NAND2_X1 U173 ( .A1(n179), .A2(n40), .ZN(n5) );
  NAND2_X1 U174 ( .A1(n94), .A2(n33), .ZN(n4) );
  NAND2_X1 U175 ( .A1(n93), .A2(n26), .ZN(n3) );
  INV_X1 U176 ( .A(n25), .ZN(n93) );
  NOR2_X1 U177 ( .A1(n163), .A2(n42), .ZN(n37) );
  XNOR2_X1 U178 ( .A(n10), .B(n65), .ZN(SUM[7]) );
  NAND2_X1 U179 ( .A1(n173), .A2(n64), .ZN(n10) );
  XNOR2_X1 U180 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U181 ( .A1(n186), .A2(n19), .ZN(n2) );
  NAND2_X1 U182 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  INV_X1 U183 ( .A(n32), .ZN(n94) );
  OAI21_X1 U184 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  NOR2_X1 U185 ( .A1(n32), .A2(n25), .ZN(n23) );
  INV_X1 U186 ( .A(n64), .ZN(n62) );
  OR2_X1 U187 ( .A1(B[15]), .A2(A[15]), .ZN(n186) );
  NOR2_X1 U188 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  XNOR2_X1 U189 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  NAND2_X1 U190 ( .A1(n189), .A2(n78), .ZN(n13) );
  NOR2_X1 U191 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  INV_X1 U192 ( .A(n80), .ZN(n104) );
  NOR2_X1 U193 ( .A1(A[12]), .A2(B[12]), .ZN(n39) );
  NAND2_X1 U194 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  OAI21_X1 U195 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  AOI21_X1 U196 ( .B1(n189), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U197 ( .A(n78), .ZN(n76) );
  OR2_X1 U198 ( .A1(B[2]), .A2(A[2]), .ZN(n187) );
  NOR2_X1 U199 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  NAND2_X1 U200 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  NAND2_X1 U201 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  OR2_X1 U202 ( .A1(B[6]), .A2(A[6]), .ZN(n188) );
  NAND2_X1 U203 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND2_X1 U204 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  XNOR2_X1 U205 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U206 ( .A1(n187), .A2(n86), .ZN(n15) );
  AOI21_X1 U207 ( .B1(n87), .B2(n187), .A(n84), .ZN(n82) );
  INV_X1 U208 ( .A(n86), .ZN(n84) );
  NOR2_X1 U209 ( .A1(B[3]), .A2(A[3]), .ZN(n80) );
  OR2_X1 U210 ( .A1(B[4]), .A2(A[4]), .ZN(n189) );
  NAND2_X1 U211 ( .A1(B[3]), .A2(A[3]), .ZN(n81) );
  XOR2_X1 U212 ( .A(n16), .B(n91), .Z(SUM[1]) );
  INV_X1 U213 ( .A(n88), .ZN(n106) );
  OAI21_X1 U214 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U215 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U216 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  NAND2_X1 U217 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  NAND2_X1 U218 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  NAND2_X1 U219 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  NAND2_X1 U220 ( .A1(n106), .A2(n89), .ZN(n16) );
  NAND2_X1 U221 ( .A1(n104), .A2(n81), .ZN(n14) );
  XOR2_X1 U222 ( .A(n14), .B(n82), .Z(SUM[3]) );
  XNOR2_X1 U223 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U224 ( .A1(n37), .A2(n94), .ZN(n28) );
  INV_X1 U225 ( .A(n37), .ZN(n35) );
  INV_X1 U226 ( .A(n38), .ZN(n36) );
  AOI21_X1 U227 ( .B1(n38), .B2(n94), .A(n31), .ZN(n29) );
  OAI21_X1 U228 ( .B1(n54), .B2(n66), .A(n55), .ZN(n53) );
  NAND2_X1 U229 ( .A1(n102), .A2(n73), .ZN(n12) );
  NAND2_X1 U230 ( .A1(A[9]), .A2(B[9]), .ZN(n51) );
  AOI21_X1 U231 ( .B1(n65), .B2(n173), .A(n62), .ZN(n60) );
  XNOR2_X1 U232 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U233 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
  NAND2_X1 U234 ( .A1(n170), .A2(n23), .ZN(n21) );
  AOI21_X1 U235 ( .B1(n23), .B2(n167), .A(n24), .ZN(n22) );
  OAI21_X1 U236 ( .B1(n178), .B2(n52), .A(n177), .ZN(n49) );
  NAND2_X1 U237 ( .A1(A[7]), .A2(B[7]), .ZN(n64) );
  INV_X1 U238 ( .A(n53), .ZN(n52) );
  NAND2_X1 U239 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  OAI21_X1 U240 ( .B1(n21), .B2(n162), .A(n22), .ZN(n20) );
  OAI21_X1 U241 ( .B1(n28), .B2(n171), .A(n29), .ZN(n27) );
  OAI21_X1 U242 ( .B1(n171), .B2(n165), .A(n43), .ZN(n41) );
  XNOR2_X1 U243 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  OAI21_X1 U244 ( .B1(n35), .B2(n1), .A(n36), .ZN(n34) );
  OAI21_X1 U245 ( .B1(n47), .B2(n51), .A(n48), .ZN(n46) );
  NOR2_X1 U246 ( .A1(n181), .A2(n178), .ZN(n45) );
  AOI21_X1 U247 ( .B1(n190), .B2(n62), .A(n176), .ZN(n55) );
  NAND2_X1 U248 ( .A1(n168), .A2(n173), .ZN(n54) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_0 ( .in({\in[3][15] , 
        \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , \in[3][10] , 
        \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , \in[3][5] , \in[3][4] , 
        \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , \in[2][15] , 
        \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , \in[2][10] , 
        \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , \in[2][5] , \in[2][4] , 
        \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , \in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \genblk1.inter[1][15] , \genblk1.inter[1][14] ,
         \genblk1.inter[1][13] , \genblk1.inter[1][12] ,
         \genblk1.inter[1][11] , \genblk1.inter[1][10] , \genblk1.inter[1][9] ,
         \genblk1.inter[1][8] , \genblk1.inter[1][7] , \genblk1.inter[1][6] ,
         \genblk1.inter[1][5] , \genblk1.inter[1][4] , \genblk1.inter[1][3] ,
         \genblk1.inter[1][2] , \genblk1.inter[1][1] , \genblk1.inter[1][0] ,
         \genblk1.inter[0][15] , \genblk1.inter[0][14] ,
         \genblk1.inter[0][13] , \genblk1.inter[0][12] ,
         \genblk1.inter[0][11] , \genblk1.inter[0][10] , \genblk1.inter[0][9] ,
         \genblk1.inter[0][8] , \genblk1.inter[0][7] , \genblk1.inter[0][6] ,
         \genblk1.inter[0][5] , \genblk1.inter[0][4] , \genblk1.inter[0][3] ,
         \genblk1.inter[0][2] , \genblk1.inter[0][1] , \genblk1.inter[0][0] ;

  recursive_add_layer_INPUT_SCALE2_WIDTH16_0 \genblk1.next_layer  ( .in({
        \genblk1.inter[1][15] , \genblk1.inter[1][14] , \genblk1.inter[1][13] , 
        \genblk1.inter[1][12] , \genblk1.inter[1][11] , \genblk1.inter[1][10] , 
        \genblk1.inter[1][9] , \genblk1.inter[1][8] , \genblk1.inter[1][7] , 
        \genblk1.inter[1][6] , \genblk1.inter[1][5] , \genblk1.inter[1][4] , 
        \genblk1.inter[1][3] , \genblk1.inter[1][2] , \genblk1.inter[1][1] , 
        \genblk1.inter[1][0] , \genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }), .out(out) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_0_DW01_add_4 add_64_G2 ( .A({
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] }), .B({\in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] }), .CI(1'b0), .SUM({\genblk1.inter[1][15] , \genblk1.inter[1][14] , 
        \genblk1.inter[1][13] , \genblk1.inter[1][12] , \genblk1.inter[1][11] , 
        \genblk1.inter[1][10] , \genblk1.inter[1][9] , \genblk1.inter[1][8] , 
        \genblk1.inter[1][7] , \genblk1.inter[1][6] , \genblk1.inter[1][5] , 
        \genblk1.inter[1][4] , \genblk1.inter[1][3] , \genblk1.inter[1][2] , 
        \genblk1.inter[1][1] , \genblk1.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_0_DW01_add_5 add_64 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM({\genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }) );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_0 ( .a({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , 
        \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , 
        \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , 
        \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , \x[1][7] , 
        \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , 
        \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , 
        \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \multout[3][15] , \multout[3][14] , \multout[3][13] ,
         \multout[3][12] , \multout[3][11] , \multout[3][10] , \multout[3][9] ,
         \multout[3][8] , \multout[3][7] , \multout[3][6] , \multout[3][5] ,
         \multout[3][4] , \multout[3][3] , \multout[3][2] , \multout[3][1] ,
         \multout[3][0] , \multout[2][15] , \multout[2][14] , \multout[2][13] ,
         \multout[2][12] , \multout[2][11] , \multout[2][10] , \multout[2][9] ,
         \multout[2][8] , \multout[2][7] , \multout[2][6] , \multout[2][5] ,
         \multout[2][4] , \multout[2][3] , \multout[2][2] , \multout[2][1] ,
         \multout[2][0] , \multout[1][15] , \multout[1][14] , \multout[1][13] ,
         \multout[1][12] , \multout[1][11] , \multout[1][10] , \multout[1][9] ,
         \multout[1][8] , \multout[1][7] , \multout[1][6] , \multout[1][5] ,
         \multout[1][4] , \multout[1][3] , \multout[1][2] , \multout[1][1] ,
         \multout[1][0] , \multout[0][15] , \multout[0][14] , \multout[0][13] ,
         \multout[0][12] , \multout[0][11] , \multout[0][10] , \multout[0][9] ,
         \multout[0][8] , \multout[0][7] , \multout[0][6] , \multout[0][5] ,
         \multout[0][4] , \multout[0][3] , \multout[0][2] , \multout[0][1] ,
         \multout[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_0 \genblk1[0].mult  ( .ia({\a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({\multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_15 \genblk1[1].mult  ( .ia({\a[1][7] , 
        \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , 
        \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , 
        \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({\multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_14 \genblk1[2].mult  ( .ia({\a[2][7] , 
        \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , \a[2][1] , 
        \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] , 
        \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({\multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_13 \genblk1[3].mult  ( .ia({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_0 add ( .in({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] , \multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] , \multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] , \multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102,
         n103, n104, n109, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n163, n164, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n245, n246, n247, n248, n250, n251, n252,
         n253, n254, n255, n256, n258, n259, n260, n261, n262, n263, n264,
         n265, n273, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n356,
         n357;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n325), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U141 ( .A(n195), .B(n182), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n199), .B(n192), .CO(n152), .S(n153) );
  XOR2_X1 U268 ( .A(b[7]), .B(n261), .Z(n229) );
  CLKBUF_X1 U269 ( .A(n265), .Z(n338) );
  CLKBUF_X1 U270 ( .A(n262), .Z(n303) );
  NOR2_X1 U271 ( .A1(n121), .A2(n124), .ZN(n304) );
  NOR2_X1 U272 ( .A1(n121), .A2(n124), .ZN(n61) );
  CLKBUF_X1 U273 ( .A(n265), .Z(n305) );
  CLKBUF_X1 U274 ( .A(n74), .Z(n306) );
  XNOR2_X1 U275 ( .A(n265), .B(n164), .ZN(n307) );
  BUF_X1 U276 ( .A(n264), .Z(n308) );
  BUF_X1 U277 ( .A(n141), .Z(n309) );
  BUF_X2 U278 ( .A(n263), .Z(n318) );
  CLKBUF_X1 U279 ( .A(n264), .Z(n310) );
  CLKBUF_X1 U280 ( .A(n354), .Z(n311) );
  CLKBUF_X1 U281 ( .A(n265), .Z(n312) );
  OR2_X1 U282 ( .A1(n151), .A2(n152), .ZN(n313) );
  CLKBUF_X1 U283 ( .A(n88), .Z(n314) );
  INV_X1 U284 ( .A(n57), .ZN(n315) );
  NOR2_X1 U285 ( .A1(n64), .A2(n61), .ZN(n3) );
  XNOR2_X1 U286 ( .A(n264), .B(a[4]), .ZN(n316) );
  OAI21_X1 U287 ( .B1(n61), .B2(n65), .A(n62), .ZN(n317) );
  OAI21_X1 U288 ( .B1(n304), .B2(n65), .A(n62), .ZN(n2) );
  XNOR2_X2 U289 ( .A(n265), .B(a[2]), .ZN(n324) );
  XNOR2_X1 U290 ( .A(n133), .B(n319), .ZN(n131) );
  XNOR2_X1 U291 ( .A(n138), .B(n135), .ZN(n319) );
  XOR2_X1 U292 ( .A(n141), .B(n144), .Z(n320) );
  XOR2_X1 U293 ( .A(n139), .B(n320), .Z(n137) );
  NAND2_X1 U294 ( .A1(n139), .A2(n144), .ZN(n321) );
  NAND2_X1 U295 ( .A1(n139), .A2(n309), .ZN(n322) );
  NAND2_X1 U296 ( .A1(n144), .A2(n141), .ZN(n323) );
  NAND3_X1 U297 ( .A1(n321), .A2(n322), .A3(n323), .ZN(n136) );
  OAI22_X1 U298 ( .A1(n344), .A2(n221), .B1(n220), .B2(n324), .ZN(n325) );
  BUF_X1 U299 ( .A(n252), .Z(n344) );
  OR2_X1 U300 ( .A1(n201), .A2(n169), .ZN(n326) );
  INV_X1 U301 ( .A(n259), .ZN(n327) );
  NAND2_X1 U302 ( .A1(n133), .A2(n138), .ZN(n328) );
  NAND2_X1 U303 ( .A1(n133), .A2(n135), .ZN(n329) );
  NAND2_X1 U304 ( .A1(n138), .A2(n135), .ZN(n330) );
  NAND3_X1 U305 ( .A1(n328), .A2(n329), .A3(n330), .ZN(n130) );
  NAND2_X1 U306 ( .A1(n246), .A2(n254), .ZN(n331) );
  XNOR2_X1 U307 ( .A(n263), .B(a[6]), .ZN(n332) );
  BUF_X1 U308 ( .A(n252), .Z(n343) );
  XOR2_X1 U309 ( .A(a[6]), .B(n262), .Z(n333) );
  CLKBUF_X1 U310 ( .A(n262), .Z(n334) );
  CLKBUF_X1 U311 ( .A(n83), .Z(n335) );
  XNOR2_X1 U312 ( .A(n356), .B(n336), .ZN(product[9]) );
  AND2_X1 U313 ( .A1(n103), .A2(n65), .ZN(n336) );
  INV_X1 U314 ( .A(n340), .ZN(n82) );
  OR2_X1 U315 ( .A1(n137), .A2(n142), .ZN(n337) );
  OR2_X2 U316 ( .A1(n307), .A2(n164), .ZN(n339) );
  XNOR2_X1 U317 ( .A(n263), .B(a[6]), .ZN(n352) );
  BUF_X2 U318 ( .A(n1), .Z(n356) );
  AND2_X1 U319 ( .A1(n147), .A2(n150), .ZN(n340) );
  FA_X1 U320 ( .A(n148), .B(n183), .CI(n145), .S(n341) );
  OR2_X1 U321 ( .A1(n341), .A2(n146), .ZN(n342) );
  NAND2_X1 U322 ( .A1(n248), .A2(n256), .ZN(n252) );
  INV_X1 U323 ( .A(n260), .ZN(n345) );
  NOR2_X1 U324 ( .A1(n131), .A2(n136), .ZN(n346) );
  NOR2_X1 U325 ( .A1(n131), .A2(n136), .ZN(n69) );
  XNOR2_X1 U326 ( .A(n264), .B(a[4]), .ZN(n347) );
  BUF_X2 U327 ( .A(n245), .Z(n357) );
  NAND2_X1 U328 ( .A1(n333), .A2(n332), .ZN(n348) );
  CLKBUF_X1 U329 ( .A(n78), .Z(n349) );
  OR2_X2 U330 ( .A1(n350), .A2(n164), .ZN(n253) );
  XNOR2_X1 U331 ( .A(n265), .B(n164), .ZN(n350) );
  INV_X1 U332 ( .A(n164), .ZN(n273) );
  NAND2_X1 U333 ( .A1(n247), .A2(n255), .ZN(n351) );
  INV_X1 U334 ( .A(n30), .ZN(n28) );
  INV_X1 U335 ( .A(n64), .ZN(n103) );
  INV_X1 U336 ( .A(n18), .ZN(product[15]) );
  AOI21_X1 U337 ( .B1(n317), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U338 ( .B1(n317), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U339 ( .A(n31), .ZN(n29) );
  INV_X1 U340 ( .A(n317), .ZN(n58) );
  NAND2_X1 U341 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U342 ( .A(n304), .ZN(n102) );
  NAND2_X1 U343 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U344 ( .A(n41), .ZN(n100) );
  NAND2_X1 U345 ( .A1(n337), .A2(n73), .ZN(n11) );
  XNOR2_X1 U346 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U347 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U348 ( .A(n34), .ZN(n99) );
  NAND2_X1 U349 ( .A1(n311), .A2(n82), .ZN(n13) );
  AOI21_X1 U350 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U351 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U352 ( .A(n56), .B(n7), .ZN(product[11]) );
  XNOR2_X1 U353 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U354 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U355 ( .A(n23), .ZN(n98) );
  NOR2_X1 U356 ( .A1(n125), .A2(n130), .ZN(n64) );
  NAND2_X1 U357 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U358 ( .A(n346), .ZN(n104) );
  AOI21_X1 U359 ( .B1(n353), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U360 ( .A(n94), .ZN(n92) );
  OAI21_X1 U361 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  OAI21_X1 U362 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  NOR2_X1 U363 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U364 ( .A1(n50), .A2(n41), .ZN(n39) );
  NOR2_X1 U365 ( .A1(n41), .A2(n34), .ZN(n32) );
  NAND2_X1 U366 ( .A1(n125), .A2(n130), .ZN(n65) );
  AOI21_X1 U367 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U368 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  INV_X1 U369 ( .A(n51), .ZN(n53) );
  NAND2_X1 U370 ( .A1(n131), .A2(n136), .ZN(n70) );
  INV_X1 U371 ( .A(n50), .ZN(n52) );
  XNOR2_X1 U372 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U373 ( .A1(n353), .A2(n94), .ZN(n16) );
  NAND2_X1 U374 ( .A1(n342), .A2(n77), .ZN(n12) );
  XOR2_X1 U375 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U376 ( .A1(n313), .A2(n85), .ZN(n14) );
  XOR2_X1 U377 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U378 ( .A(n314), .ZN(n109) );
  NOR2_X1 U379 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U380 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U381 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U382 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U383 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U384 ( .A(n112), .ZN(n113) );
  NOR2_X1 U385 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U386 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U387 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U388 ( .A1(n137), .A2(n142), .ZN(n72) );
  INV_X1 U389 ( .A(n97), .ZN(n95) );
  OR2_X1 U390 ( .A1(n200), .A2(n193), .ZN(n353) );
  NOR2_X1 U391 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U392 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U393 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U394 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U395 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U396 ( .A1(n341), .A2(n146), .ZN(n77) );
  OR2_X1 U397 ( .A1(n147), .A2(n150), .ZN(n354) );
  INV_X1 U398 ( .A(n87), .ZN(n86) );
  AND2_X1 U399 ( .A1(n357), .A2(n161), .ZN(n193) );
  INV_X1 U400 ( .A(n157), .ZN(n178) );
  OAI22_X1 U401 ( .A1(n339), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  AND2_X1 U402 ( .A1(n357), .A2(n158), .ZN(n185) );
  OAI22_X1 U403 ( .A1(n339), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  INV_X1 U404 ( .A(n118), .ZN(n119) );
  OR2_X1 U405 ( .A1(n357), .A2(n259), .ZN(n219) );
  AND2_X1 U406 ( .A1(n326), .A2(n97), .ZN(product[1]) );
  INV_X1 U407 ( .A(n163), .ZN(n194) );
  OAI22_X1 U408 ( .A1(n339), .A2(n229), .B1(n229), .B2(n273), .ZN(n163) );
  INV_X1 U409 ( .A(n160), .ZN(n186) );
  INV_X1 U410 ( .A(n128), .ZN(n129) );
  OAI22_X1 U411 ( .A1(n339), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  AND2_X1 U412 ( .A1(n357), .A2(n155), .ZN(n177) );
  OAI22_X1 U413 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  NOR2_X1 U414 ( .A1(n151), .A2(n152), .ZN(n84) );
  NOR2_X1 U415 ( .A1(n153), .A2(n168), .ZN(n88) );
  INV_X1 U416 ( .A(n154), .ZN(n170) );
  NAND2_X1 U417 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U418 ( .A1(n357), .A2(n258), .ZN(n210) );
  XNOR2_X1 U419 ( .A(n263), .B(a[6]), .ZN(n254) );
  OR2_X1 U420 ( .A1(n357), .A2(n260), .ZN(n228) );
  OAI22_X1 U421 ( .A1(n339), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OR2_X1 U422 ( .A1(n357), .A2(n261), .ZN(n237) );
  OAI22_X1 U423 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  XNOR2_X1 U424 ( .A(b[7]), .B(n334), .ZN(n202) );
  NAND2_X1 U425 ( .A1(n246), .A2(n254), .ZN(n250) );
  XOR2_X1 U426 ( .A(a[6]), .B(n262), .Z(n246) );
  XNOR2_X1 U427 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U428 ( .A(b[4]), .B(n303), .ZN(n205) );
  XNOR2_X1 U429 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U430 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U431 ( .A(b[6]), .B(n262), .ZN(n203) );
  NAND2_X1 U432 ( .A1(n247), .A2(n255), .ZN(n251) );
  XNOR2_X1 U433 ( .A(b[1]), .B(n262), .ZN(n208) );
  AND2_X1 U434 ( .A1(n357), .A2(n164), .ZN(product[0]) );
  XNOR2_X1 U435 ( .A(n262), .B(n357), .ZN(n209) );
  INV_X1 U436 ( .A(n262), .ZN(n258) );
  AOI21_X1 U437 ( .B1(n75), .B2(n67), .A(n68), .ZN(n1) );
  NAND2_X1 U438 ( .A1(n200), .A2(n193), .ZN(n94) );
  OAI22_X1 U439 ( .A1(n339), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  XNOR2_X1 U440 ( .A(n264), .B(a[4]), .ZN(n255) );
  NAND2_X1 U441 ( .A1(n315), .A2(n21), .ZN(n19) );
  NAND2_X1 U442 ( .A1(n315), .A2(n28), .ZN(n26) );
  NAND2_X1 U443 ( .A1(n3), .A2(n39), .ZN(n37) );
  INV_X1 U444 ( .A(n3), .ZN(n57) );
  OAI21_X1 U445 ( .B1(n356), .B2(n19), .A(n20), .ZN(n18) );
  XNOR2_X1 U446 ( .A(n63), .B(n8), .ZN(product[10]) );
  NOR2_X1 U447 ( .A1(n346), .A2(n72), .ZN(n67) );
  NAND2_X1 U448 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U449 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  XNOR2_X1 U450 ( .A(n71), .B(n10), .ZN(product[8]) );
  XNOR2_X1 U451 ( .A(n13), .B(n335), .ZN(product[5]) );
  AOI21_X1 U452 ( .B1(n354), .B2(n83), .A(n340), .ZN(n78) );
  OAI21_X1 U453 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  OAI21_X1 U454 ( .B1(n64), .B2(n1), .A(n65), .ZN(n63) );
  OAI21_X1 U455 ( .B1(n356), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U456 ( .B1(n356), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U457 ( .B1(n356), .B2(n26), .A(n27), .ZN(n25) );
  NAND2_X1 U458 ( .A1(n52), .A2(n51), .ZN(n7) );
  NAND2_X1 U459 ( .A1(n3), .A2(n52), .ZN(n46) );
  AOI21_X1 U460 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  NAND2_X1 U461 ( .A1(n52), .A2(n32), .ZN(n30) );
  XOR2_X1 U462 ( .A(n306), .B(n11), .Z(product[7]) );
  OAI21_X1 U463 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  INV_X1 U464 ( .A(n75), .ZN(n74) );
  OAI21_X1 U465 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NAND2_X1 U466 ( .A1(n109), .A2(n89), .ZN(n15) );
  XNOR2_X1 U467 ( .A(n45), .B(n6), .ZN(product[12]) );
  OAI21_X1 U468 ( .B1(n46), .B2(n356), .A(n47), .ZN(n45) );
  OAI21_X1 U469 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  OAI22_X1 U470 ( .A1(n343), .A2(n225), .B1(n224), .B2(n324), .ZN(n190) );
  OAI22_X1 U471 ( .A1(n343), .A2(n260), .B1(n228), .B2(n324), .ZN(n168) );
  OAI22_X1 U472 ( .A1(n343), .A2(n222), .B1(n221), .B2(n324), .ZN(n187) );
  OAI22_X1 U473 ( .A1(n252), .A2(n224), .B1(n324), .B2(n223), .ZN(n189) );
  OAI22_X1 U474 ( .A1(n343), .A2(n223), .B1(n222), .B2(n324), .ZN(n188) );
  OAI22_X1 U475 ( .A1(n344), .A2(n226), .B1(n225), .B2(n324), .ZN(n191) );
  OAI22_X1 U476 ( .A1(n343), .A2(n221), .B1(n220), .B2(n324), .ZN(n128) );
  OAI22_X1 U477 ( .A1(n220), .A2(n344), .B1(n220), .B2(n324), .ZN(n160) );
  XNOR2_X1 U478 ( .A(b[5]), .B(n265), .ZN(n231) );
  XNOR2_X1 U479 ( .A(n265), .B(b[6]), .ZN(n230) );
  XNOR2_X1 U480 ( .A(b[4]), .B(n338), .ZN(n232) );
  OAI22_X1 U481 ( .A1(n252), .A2(n227), .B1(n226), .B2(n324), .ZN(n192) );
  INV_X1 U482 ( .A(n324), .ZN(n161) );
  XNOR2_X1 U483 ( .A(b[3]), .B(n305), .ZN(n233) );
  XNOR2_X1 U484 ( .A(n338), .B(n357), .ZN(n236) );
  XNOR2_X1 U485 ( .A(b[2]), .B(n338), .ZN(n234) );
  XNOR2_X1 U486 ( .A(b[1]), .B(n312), .ZN(n235) );
  INV_X1 U487 ( .A(n265), .ZN(n261) );
  XNOR2_X1 U488 ( .A(n265), .B(a[2]), .ZN(n256) );
  OAI22_X1 U489 ( .A1(n351), .A2(n217), .B1(n216), .B2(n347), .ZN(n183) );
  OAI22_X1 U490 ( .A1(n351), .A2(n212), .B1(n211), .B2(n347), .ZN(n118) );
  OAI22_X1 U491 ( .A1(n211), .A2(n351), .B1(n211), .B2(n316), .ZN(n157) );
  OAI22_X1 U492 ( .A1(n351), .A2(n213), .B1(n212), .B2(n347), .ZN(n179) );
  OAI22_X1 U493 ( .A1(n351), .A2(n214), .B1(n213), .B2(n347), .ZN(n180) );
  OAI22_X1 U494 ( .A1(n351), .A2(n216), .B1(n215), .B2(n347), .ZN(n182) );
  OAI22_X1 U495 ( .A1(n351), .A2(n215), .B1(n214), .B2(n316), .ZN(n181) );
  INV_X1 U496 ( .A(n347), .ZN(n158) );
  OAI22_X1 U497 ( .A1(n251), .A2(n259), .B1(n219), .B2(n316), .ZN(n167) );
  OAI22_X1 U498 ( .A1(n251), .A2(n218), .B1(n217), .B2(n316), .ZN(n184) );
  XNOR2_X1 U499 ( .A(b[3]), .B(n308), .ZN(n224) );
  XNOR2_X1 U500 ( .A(b[5]), .B(n310), .ZN(n222) );
  XNOR2_X1 U501 ( .A(b[4]), .B(n308), .ZN(n223) );
  INV_X1 U502 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U503 ( .A(b[2]), .B(n345), .ZN(n225) );
  XNOR2_X1 U504 ( .A(b[6]), .B(n345), .ZN(n221) );
  XNOR2_X1 U505 ( .A(b[7]), .B(n310), .ZN(n220) );
  XNOR2_X1 U506 ( .A(n345), .B(n357), .ZN(n227) );
  XNOR2_X1 U507 ( .A(b[1]), .B(n308), .ZN(n226) );
  XOR2_X1 U508 ( .A(n264), .B(a[2]), .Z(n248) );
  OAI22_X1 U509 ( .A1(n202), .A2(n331), .B1(n202), .B2(n254), .ZN(n154) );
  OAI22_X1 U510 ( .A1(n331), .A2(n206), .B1(n205), .B2(n332), .ZN(n173) );
  OAI22_X1 U511 ( .A1(n348), .A2(n203), .B1(n202), .B2(n332), .ZN(n112) );
  OAI22_X1 U512 ( .A1(n331), .A2(n205), .B1(n204), .B2(n254), .ZN(n172) );
  OAI22_X1 U513 ( .A1(n348), .A2(n204), .B1(n203), .B2(n254), .ZN(n171) );
  OAI22_X1 U514 ( .A1(n348), .A2(n207), .B1(n206), .B2(n352), .ZN(n174) );
  XNOR2_X1 U515 ( .A(b[7]), .B(n327), .ZN(n211) );
  XNOR2_X1 U516 ( .A(b[6]), .B(n327), .ZN(n212) );
  INV_X1 U517 ( .A(n352), .ZN(n155) );
  XNOR2_X1 U518 ( .A(b[5]), .B(n318), .ZN(n213) );
  OAI22_X1 U519 ( .A1(n331), .A2(n208), .B1(n207), .B2(n352), .ZN(n175) );
  OAI22_X1 U520 ( .A1(n348), .A2(n258), .B1(n352), .B2(n210), .ZN(n166) );
  OAI22_X1 U521 ( .A1(n250), .A2(n209), .B1(n208), .B2(n352), .ZN(n176) );
  XNOR2_X1 U522 ( .A(b[2]), .B(n318), .ZN(n216) );
  XNOR2_X1 U523 ( .A(b[3]), .B(n318), .ZN(n215) );
  XNOR2_X1 U524 ( .A(b[4]), .B(n327), .ZN(n214) );
  XNOR2_X1 U525 ( .A(n318), .B(n357), .ZN(n218) );
  INV_X1 U526 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U527 ( .A(b[1]), .B(n318), .ZN(n217) );
  XOR2_X1 U528 ( .A(n263), .B(a[4]), .Z(n247) );
  XOR2_X1 U529 ( .A(n12), .B(n349), .Z(product[6]) );
  NAND2_X1 U530 ( .A1(n153), .A2(n168), .ZN(n89) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n12, n13, n14, n15, n16, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50,
         n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102, n103,
         n104, n105, n106, n109, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n157, n158, n160, n161, n163, n164, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n245, n246, n247, n248, n250, n251, n252,
         n253, n254, n255, n256, n258, n259, n260, n261, n262, n263, n264,
         n265, n273, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n370, n371, n372;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U136 ( .A(n138), .B(n135), .CI(n133), .CO(n130), .S(n131) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U144 ( .A(n177), .B(n189), .CI(n196), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n199), .B(n192), .CO(n152), .S(n153) );
  XNOR2_X1 U268 ( .A(n264), .B(a[4]), .ZN(n303) );
  BUF_X1 U269 ( .A(n341), .Z(n304) );
  CLKBUF_X2 U270 ( .A(n263), .Z(n350) );
  XOR2_X1 U271 ( .A(n179), .B(n341), .Z(n305) );
  XOR2_X1 U272 ( .A(n305), .B(n186), .Z(n123) );
  XOR2_X1 U273 ( .A(n126), .B(n173), .Z(n306) );
  XOR2_X1 U274 ( .A(n306), .B(n123), .Z(n121) );
  NAND2_X1 U275 ( .A1(n179), .A2(n304), .ZN(n307) );
  NAND2_X1 U276 ( .A1(n179), .A2(n186), .ZN(n308) );
  NAND2_X1 U277 ( .A1(n304), .A2(n186), .ZN(n309) );
  NAND3_X1 U278 ( .A1(n307), .A2(n308), .A3(n309), .ZN(n122) );
  NAND2_X1 U279 ( .A1(n126), .A2(n173), .ZN(n310) );
  NAND2_X1 U280 ( .A1(n126), .A2(n123), .ZN(n311) );
  NAND2_X1 U281 ( .A1(n173), .A2(n123), .ZN(n312) );
  NAND3_X1 U282 ( .A1(n310), .A2(n311), .A3(n312), .ZN(n120) );
  CLKBUF_X1 U283 ( .A(n264), .Z(n313) );
  CLKBUF_X1 U284 ( .A(n371), .Z(n314) );
  OR2_X1 U285 ( .A1(n151), .A2(n152), .ZN(n315) );
  NAND2_X2 U286 ( .A1(n248), .A2(n256), .ZN(n364) );
  OR2_X1 U287 ( .A1(n147), .A2(n150), .ZN(n316) );
  INV_X1 U288 ( .A(n335), .ZN(n317) );
  CLKBUF_X1 U289 ( .A(n313), .Z(n318) );
  NAND2_X1 U290 ( .A1(n337), .A2(n338), .ZN(n319) );
  CLKBUF_X1 U291 ( .A(n344), .Z(n320) );
  CLKBUF_X1 U292 ( .A(n262), .Z(n321) );
  XOR2_X1 U293 ( .A(n199), .B(n192), .Z(n322) );
  OAI22_X2 U294 ( .A1(n252), .A2(n227), .B1(n226), .B2(n333), .ZN(n192) );
  INV_X1 U295 ( .A(n259), .ZN(n323) );
  XOR2_X1 U296 ( .A(n144), .B(n141), .Z(n324) );
  XOR2_X1 U297 ( .A(n139), .B(n324), .Z(n137) );
  NAND2_X1 U298 ( .A1(n139), .A2(n144), .ZN(n325) );
  NAND2_X1 U299 ( .A1(n139), .A2(n141), .ZN(n326) );
  NAND2_X1 U300 ( .A1(n144), .A2(n141), .ZN(n327) );
  NAND3_X1 U301 ( .A1(n325), .A2(n326), .A3(n327), .ZN(n136) );
  XNOR2_X2 U302 ( .A(n263), .B(a[6]), .ZN(n366) );
  XOR2_X1 U303 ( .A(n148), .B(n183), .Z(n328) );
  XOR2_X1 U304 ( .A(n145), .B(n328), .Z(n143) );
  NAND2_X1 U305 ( .A1(n145), .A2(n148), .ZN(n329) );
  NAND2_X1 U306 ( .A1(n145), .A2(n183), .ZN(n330) );
  NAND2_X1 U307 ( .A1(n148), .A2(n183), .ZN(n331) );
  NAND3_X1 U308 ( .A1(n329), .A2(n330), .A3(n331), .ZN(n142) );
  AND2_X1 U309 ( .A1(n147), .A2(n150), .ZN(n332) );
  XNOR2_X1 U310 ( .A(n265), .B(a[2]), .ZN(n333) );
  CLKBUF_X1 U311 ( .A(n264), .Z(n334) );
  NOR2_X1 U312 ( .A1(n347), .A2(n72), .ZN(n67) );
  NAND2_X1 U313 ( .A1(a[6]), .A2(n336), .ZN(n337) );
  NAND2_X1 U314 ( .A1(n335), .A2(n262), .ZN(n338) );
  NAND2_X1 U315 ( .A1(n337), .A2(n338), .ZN(n246) );
  INV_X1 U316 ( .A(a[6]), .ZN(n335) );
  INV_X1 U317 ( .A(n262), .ZN(n336) );
  NOR2_X1 U318 ( .A1(n64), .A2(n61), .ZN(n339) );
  BUF_X1 U319 ( .A(n362), .Z(n340) );
  NOR2_X2 U320 ( .A1(n121), .A2(n124), .ZN(n61) );
  OAI22_X1 U321 ( .A1(n364), .A2(n221), .B1(n220), .B2(n333), .ZN(n341) );
  OAI21_X1 U322 ( .B1(n61), .B2(n65), .A(n62), .ZN(n342) );
  BUF_X2 U323 ( .A(n245), .Z(n372) );
  OAI21_X1 U324 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  OR2_X1 U325 ( .A1(n201), .A2(n169), .ZN(n343) );
  AND2_X1 U326 ( .A1(n105), .A2(n73), .ZN(n351) );
  AOI21_X1 U327 ( .B1(n67), .B2(n363), .A(n68), .ZN(n344) );
  AOI21_X1 U328 ( .B1(n67), .B2(n363), .A(n68), .ZN(n345) );
  AOI21_X1 U329 ( .B1(n67), .B2(n363), .A(n68), .ZN(n365) );
  CLKBUF_X1 U330 ( .A(n265), .Z(n346) );
  NOR2_X1 U331 ( .A1(n131), .A2(n136), .ZN(n347) );
  NOR2_X1 U332 ( .A1(n131), .A2(n136), .ZN(n69) );
  OR2_X2 U333 ( .A1(n348), .A2(n164), .ZN(n253) );
  XNOR2_X1 U334 ( .A(n265), .B(n164), .ZN(n348) );
  INV_X1 U335 ( .A(n164), .ZN(n273) );
  CLKBUF_X1 U336 ( .A(n83), .Z(n349) );
  OAI21_X1 U337 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  XNOR2_X1 U338 ( .A(n351), .B(n74), .ZN(product[7]) );
  NAND2_X1 U339 ( .A1(n319), .A2(n366), .ZN(n352) );
  NAND2_X1 U340 ( .A1(n319), .A2(n366), .ZN(n353) );
  NAND2_X1 U341 ( .A1(n246), .A2(n254), .ZN(n250) );
  XNOR2_X1 U342 ( .A(n344), .B(n354), .ZN(product[9]) );
  AND2_X1 U343 ( .A1(n103), .A2(n65), .ZN(n354) );
  INV_X1 U344 ( .A(n260), .ZN(n355) );
  INV_X1 U345 ( .A(n265), .ZN(n356) );
  INV_X2 U346 ( .A(n356), .ZN(n357) );
  XNOR2_X1 U347 ( .A(n264), .B(a[4]), .ZN(n362) );
  XOR2_X1 U348 ( .A(n323), .B(n317), .Z(n358) );
  OAI21_X1 U349 ( .B1(n347), .B2(n73), .A(n70), .ZN(n359) );
  CLKBUF_X1 U350 ( .A(n321), .Z(n360) );
  AOI21_X1 U351 ( .B1(n316), .B2(n83), .A(n332), .ZN(n361) );
  XNOR2_X1 U352 ( .A(n264), .B(a[4]), .ZN(n255) );
  OAI21_X1 U353 ( .B1(n76), .B2(n361), .A(n77), .ZN(n363) );
  AOI21_X1 U354 ( .B1(n67), .B2(n363), .A(n359), .ZN(n1) );
  NOR2_X1 U355 ( .A1(n64), .A2(n61), .ZN(n3) );
  INV_X1 U356 ( .A(n30), .ZN(n28) );
  INV_X1 U357 ( .A(n64), .ZN(n103) );
  INV_X1 U358 ( .A(n18), .ZN(product[15]) );
  AOI21_X1 U359 ( .B1(n342), .B2(n21), .A(n22), .ZN(n20) );
  NAND2_X1 U360 ( .A1(n339), .A2(n21), .ZN(n19) );
  AOI21_X1 U361 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  AOI21_X1 U362 ( .B1(n342), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U363 ( .A(n31), .ZN(n29) );
  NAND2_X1 U364 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U365 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U366 ( .A1(n339), .A2(n39), .ZN(n37) );
  NAND2_X1 U367 ( .A1(n339), .A2(n28), .ZN(n26) );
  INV_X1 U368 ( .A(n342), .ZN(n58) );
  XNOR2_X1 U369 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U370 ( .A1(n367), .A2(n94), .ZN(n16) );
  NAND2_X1 U371 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U372 ( .A(n41), .ZN(n100) );
  NAND2_X1 U373 ( .A1(n52), .A2(n51), .ZN(n7) );
  INV_X1 U374 ( .A(n3), .ZN(n57) );
  AOI21_X1 U375 ( .B1(n367), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U376 ( .A(n94), .ZN(n92) );
  INV_X1 U377 ( .A(n50), .ZN(n52) );
  INV_X1 U378 ( .A(n72), .ZN(n105) );
  XNOR2_X1 U379 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U380 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U381 ( .A(n23), .ZN(n98) );
  XNOR2_X1 U382 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U383 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U384 ( .A(n34), .ZN(n99) );
  NAND2_X1 U385 ( .A1(n316), .A2(n82), .ZN(n13) );
  NAND2_X1 U386 ( .A1(n104), .A2(n70), .ZN(n10) );
  AOI21_X1 U387 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U388 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  OAI21_X1 U389 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  NOR2_X1 U390 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U391 ( .A1(n125), .A2(n130), .ZN(n64) );
  NOR2_X1 U392 ( .A1(n50), .A2(n41), .ZN(n39) );
  NOR2_X1 U393 ( .A1(n41), .A2(n34), .ZN(n32) );
  NAND2_X1 U394 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U395 ( .A(n61), .ZN(n102) );
  OAI21_X1 U396 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U397 ( .A(n51), .ZN(n53) );
  NAND2_X1 U398 ( .A1(n125), .A2(n130), .ZN(n65) );
  AOI21_X1 U399 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U400 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  NAND2_X1 U401 ( .A1(n106), .A2(n77), .ZN(n12) );
  INV_X1 U402 ( .A(n76), .ZN(n106) );
  INV_X1 U403 ( .A(n88), .ZN(n109) );
  XOR2_X1 U404 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U405 ( .A1(n315), .A2(n85), .ZN(n14) );
  NOR2_X1 U406 ( .A1(n116), .A2(n115), .ZN(n41) );
  OR2_X1 U407 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U408 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U409 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U410 ( .A(n112), .ZN(n113) );
  NOR2_X1 U411 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U412 ( .A1(n170), .A2(n112), .ZN(n24) );
  XNOR2_X1 U413 ( .A(n187), .B(n175), .ZN(n135) );
  NAND2_X1 U414 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U415 ( .A1(n137), .A2(n142), .ZN(n72) );
  OAI21_X1 U416 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NOR2_X1 U417 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U418 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U419 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U420 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U421 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U422 ( .A1(n143), .A2(n146), .ZN(n77) );
  OR2_X1 U423 ( .A1(n200), .A2(n193), .ZN(n367) );
  OR2_X1 U424 ( .A1(n147), .A2(n150), .ZN(n368) );
  AND2_X1 U425 ( .A1(n372), .A2(n161), .ZN(n193) );
  INV_X1 U426 ( .A(n157), .ZN(n178) );
  INV_X1 U427 ( .A(n118), .ZN(n119) );
  AND2_X1 U428 ( .A1(n372), .A2(n158), .ZN(n185) );
  OAI22_X1 U429 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U430 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OR2_X1 U431 ( .A1(n372), .A2(n259), .ZN(n219) );
  OAI22_X1 U432 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  OAI22_X1 U433 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  INV_X1 U434 ( .A(n160), .ZN(n186) );
  INV_X1 U435 ( .A(n128), .ZN(n129) );
  OAI22_X1 U436 ( .A1(n230), .A2(n253), .B1(n229), .B2(n273), .ZN(n195) );
  AND2_X1 U437 ( .A1(n372), .A2(n358), .ZN(n177) );
  OAI22_X1 U438 ( .A1(n231), .A2(n253), .B1(n230), .B2(n273), .ZN(n196) );
  NOR2_X1 U439 ( .A1(n151), .A2(n152), .ZN(n84) );
  NAND2_X1 U440 ( .A1(n153), .A2(n168), .ZN(n89) );
  INV_X1 U441 ( .A(n154), .ZN(n170) );
  NAND2_X1 U442 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U443 ( .A1(n372), .A2(n258), .ZN(n210) );
  AND2_X1 U444 ( .A1(n343), .A2(n97), .ZN(product[1]) );
  XNOR2_X1 U445 ( .A(n263), .B(a[6]), .ZN(n254) );
  OR2_X1 U446 ( .A1(n372), .A2(n260), .ZN(n228) );
  OAI22_X1 U447 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OR2_X1 U448 ( .A1(n372), .A2(n261), .ZN(n237) );
  OAI22_X1 U449 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  XNOR2_X1 U450 ( .A(b[7]), .B(n360), .ZN(n202) );
  XNOR2_X1 U451 ( .A(b[4]), .B(n360), .ZN(n205) );
  XNOR2_X1 U452 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U453 ( .A(b[5]), .B(n360), .ZN(n204) );
  XNOR2_X1 U454 ( .A(b[6]), .B(n360), .ZN(n203) );
  NAND2_X1 U455 ( .A1(n248), .A2(n256), .ZN(n252) );
  XNOR2_X1 U456 ( .A(n262), .B(n372), .ZN(n209) );
  INV_X1 U457 ( .A(n262), .ZN(n258) );
  AND2_X1 U458 ( .A1(n372), .A2(n164), .ZN(product[0]) );
  BUF_X1 U459 ( .A(n256), .Z(n370) );
  XNOR2_X1 U460 ( .A(n265), .B(a[2]), .ZN(n256) );
  NOR2_X1 U461 ( .A1(n322), .A2(n168), .ZN(n88) );
  NAND2_X1 U462 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U463 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OAI21_X1 U464 ( .B1(n19), .B2(n320), .A(n20), .ZN(n18) );
  OAI21_X1 U465 ( .B1(n345), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U466 ( .B1(n345), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U467 ( .B1(n365), .B2(n46), .A(n47), .ZN(n45) );
  INV_X1 U468 ( .A(n163), .ZN(n194) );
  XOR2_X1 U469 ( .A(n15), .B(n90), .Z(product[3]) );
  NAND2_X1 U470 ( .A1(n109), .A2(n89), .ZN(n15) );
  INV_X1 U471 ( .A(n75), .ZN(n74) );
  INV_X1 U472 ( .A(n97), .ZN(n95) );
  XNOR2_X1 U473 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U474 ( .A1(n131), .A2(n136), .ZN(n70) );
  NAND2_X1 U475 ( .A1(n247), .A2(n362), .ZN(n371) );
  NAND2_X1 U476 ( .A1(n247), .A2(n255), .ZN(n251) );
  XNOR2_X1 U477 ( .A(n56), .B(n7), .ZN(product[11]) );
  OAI21_X1 U478 ( .B1(n365), .B2(n57), .A(n58), .ZN(n56) );
  AOI21_X1 U479 ( .B1(n368), .B2(n83), .A(n332), .ZN(n78) );
  XNOR2_X1 U480 ( .A(n13), .B(n349), .ZN(product[5]) );
  NAND2_X1 U481 ( .A1(n147), .A2(n150), .ZN(n82) );
  XNOR2_X1 U482 ( .A(n71), .B(n10), .ZN(product[8]) );
  INV_X1 U483 ( .A(n87), .ZN(n86) );
  XNOR2_X1 U484 ( .A(b[2]), .B(n321), .ZN(n207) );
  XOR2_X1 U485 ( .A(n12), .B(n361), .Z(product[6]) );
  XNOR2_X1 U486 ( .A(n63), .B(n8), .ZN(product[10]) );
  OAI21_X1 U487 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  NAND2_X1 U488 ( .A1(n200), .A2(n193), .ZN(n94) );
  XNOR2_X1 U489 ( .A(b[1]), .B(n262), .ZN(n208) );
  INV_X1 U490 ( .A(n69), .ZN(n104) );
  OAI22_X1 U491 ( .A1(n364), .A2(n260), .B1(n228), .B2(n370), .ZN(n168) );
  OAI22_X1 U492 ( .A1(n364), .A2(n222), .B1(n221), .B2(n370), .ZN(n187) );
  OAI22_X1 U493 ( .A1(n364), .A2(n225), .B1(n224), .B2(n333), .ZN(n190) );
  OAI22_X1 U494 ( .A1(n252), .A2(n224), .B1(n223), .B2(n333), .ZN(n189) );
  OAI22_X1 U495 ( .A1(n364), .A2(n226), .B1(n225), .B2(n333), .ZN(n191) );
  OAI22_X1 U496 ( .A1(n364), .A2(n221), .B1(n220), .B2(n333), .ZN(n128) );
  OAI22_X1 U497 ( .A1(n364), .A2(n223), .B1(n222), .B2(n333), .ZN(n188) );
  OAI22_X1 U498 ( .A1(n220), .A2(n364), .B1(n220), .B2(n370), .ZN(n160) );
  XNOR2_X1 U499 ( .A(b[5]), .B(n357), .ZN(n231) );
  XNOR2_X1 U500 ( .A(b[4]), .B(n357), .ZN(n232) );
  XNOR2_X1 U501 ( .A(b[6]), .B(n357), .ZN(n230) );
  INV_X1 U502 ( .A(n370), .ZN(n161) );
  XNOR2_X1 U503 ( .A(b[3]), .B(n346), .ZN(n233) );
  XNOR2_X1 U504 ( .A(n357), .B(n372), .ZN(n236) );
  XNOR2_X1 U505 ( .A(b[2]), .B(n357), .ZN(n234) );
  XNOR2_X1 U506 ( .A(b[1]), .B(n265), .ZN(n235) );
  INV_X1 U507 ( .A(n265), .ZN(n261) );
  XNOR2_X1 U508 ( .A(b[7]), .B(n346), .ZN(n229) );
  OAI21_X1 U509 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  OAI22_X1 U510 ( .A1(n371), .A2(n217), .B1(n216), .B2(n303), .ZN(n183) );
  OAI22_X1 U511 ( .A1(n314), .A2(n212), .B1(n211), .B2(n303), .ZN(n118) );
  OAI22_X1 U512 ( .A1(n211), .A2(n314), .B1(n211), .B2(n303), .ZN(n157) );
  OAI22_X1 U513 ( .A1(n371), .A2(n213), .B1(n212), .B2(n303), .ZN(n179) );
  OAI22_X1 U514 ( .A1(n371), .A2(n214), .B1(n213), .B2(n303), .ZN(n180) );
  OAI22_X1 U515 ( .A1(n371), .A2(n216), .B1(n215), .B2(n303), .ZN(n182) );
  INV_X1 U516 ( .A(n340), .ZN(n158) );
  OAI22_X1 U517 ( .A1(n371), .A2(n215), .B1(n214), .B2(n303), .ZN(n181) );
  INV_X1 U518 ( .A(n264), .ZN(n260) );
  OAI22_X1 U519 ( .A1(n251), .A2(n259), .B1(n219), .B2(n362), .ZN(n167) );
  XNOR2_X1 U520 ( .A(b[4]), .B(n264), .ZN(n223) );
  OAI22_X1 U521 ( .A1(n251), .A2(n218), .B1(n217), .B2(n340), .ZN(n184) );
  XNOR2_X1 U522 ( .A(b[3]), .B(n313), .ZN(n224) );
  XNOR2_X1 U523 ( .A(b[5]), .B(n318), .ZN(n222) );
  XNOR2_X1 U524 ( .A(b[2]), .B(n355), .ZN(n225) );
  XNOR2_X1 U525 ( .A(b[6]), .B(n355), .ZN(n221) );
  XNOR2_X1 U526 ( .A(b[7]), .B(n334), .ZN(n220) );
  XNOR2_X1 U527 ( .A(n264), .B(n372), .ZN(n227) );
  XNOR2_X1 U528 ( .A(b[1]), .B(n264), .ZN(n226) );
  XOR2_X1 U529 ( .A(n264), .B(a[2]), .Z(n248) );
  OAI22_X1 U530 ( .A1(n202), .A2(n352), .B1(n202), .B2(n366), .ZN(n154) );
  OAI22_X1 U531 ( .A1(n352), .A2(n206), .B1(n205), .B2(n366), .ZN(n173) );
  OAI22_X1 U532 ( .A1(n353), .A2(n203), .B1(n202), .B2(n366), .ZN(n112) );
  OAI22_X1 U533 ( .A1(n352), .A2(n205), .B1(n204), .B2(n366), .ZN(n172) );
  OAI22_X1 U534 ( .A1(n353), .A2(n204), .B1(n203), .B2(n366), .ZN(n171) );
  OAI22_X1 U535 ( .A1(n352), .A2(n207), .B1(n206), .B2(n366), .ZN(n174) );
  OAI22_X1 U536 ( .A1(n353), .A2(n208), .B1(n207), .B2(n366), .ZN(n175) );
  XNOR2_X1 U537 ( .A(b[7]), .B(n350), .ZN(n211) );
  XNOR2_X1 U538 ( .A(b[6]), .B(n350), .ZN(n212) );
  XNOR2_X1 U539 ( .A(b[5]), .B(n350), .ZN(n213) );
  OAI22_X1 U540 ( .A1(n250), .A2(n258), .B1(n210), .B2(n254), .ZN(n166) );
  OAI22_X1 U541 ( .A1(n250), .A2(n209), .B1(n208), .B2(n366), .ZN(n176) );
  XNOR2_X1 U542 ( .A(b[2]), .B(n350), .ZN(n216) );
  XNOR2_X1 U543 ( .A(b[3]), .B(n350), .ZN(n215) );
  XNOR2_X1 U544 ( .A(b[4]), .B(n350), .ZN(n214) );
  XNOR2_X1 U545 ( .A(n323), .B(n372), .ZN(n218) );
  INV_X1 U546 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U547 ( .A(b[1]), .B(n263), .ZN(n217) );
  XOR2_X1 U548 ( .A(n263), .B(a[4]), .Z(n247) );
  OAI21_X1 U549 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68,
         n69, n70, n71, n72, n73, n75, n76, n77, n78, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n103, n104,
         n105, n106, n108, n109, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n163, n164, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n245, n246, n247, n248, n250, n251, n253,
         n254, n255, n256, n258, n260, n261, n262, n263, n264, n265, n273,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n328), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n188), .B(n195), .CI(n182), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  CLKBUF_X1 U268 ( .A(n184), .Z(n303) );
  XNOR2_X1 U269 ( .A(n357), .B(a[4]), .ZN(n304) );
  BUF_X2 U270 ( .A(n264), .Z(n357) );
  BUF_X2 U271 ( .A(n358), .Z(n305) );
  CLKBUF_X1 U272 ( .A(n327), .Z(n306) );
  CLKBUF_X1 U273 ( .A(n65), .Z(n307) );
  NOR2_X2 U274 ( .A1(n137), .A2(n142), .ZN(n72) );
  BUF_X1 U275 ( .A(n88), .Z(n330) );
  BUF_X1 U276 ( .A(n263), .Z(n331) );
  BUF_X1 U277 ( .A(n263), .Z(n347) );
  OR2_X1 U278 ( .A1(n147), .A2(n150), .ZN(n308) );
  OR2_X1 U279 ( .A1(n147), .A2(n150), .ZN(n353) );
  OR2_X2 U280 ( .A1(n309), .A2(n164), .ZN(n253) );
  XNOR2_X1 U281 ( .A(n320), .B(n164), .ZN(n309) );
  BUF_X1 U282 ( .A(n265), .Z(n318) );
  BUF_X1 U283 ( .A(n351), .Z(n349) );
  NOR2_X1 U284 ( .A1(n121), .A2(n124), .ZN(n310) );
  NOR2_X1 U285 ( .A1(n121), .A2(n124), .ZN(n61) );
  INV_X1 U286 ( .A(n158), .ZN(n340) );
  XNOR2_X1 U287 ( .A(n306), .B(n11), .ZN(product[7]) );
  CLKBUF_X1 U288 ( .A(n265), .Z(n319) );
  CLKBUF_X1 U289 ( .A(n251), .Z(n311) );
  CLKBUF_X1 U290 ( .A(n73), .Z(n312) );
  BUF_X2 U291 ( .A(n256), .Z(n356) );
  AND2_X1 U292 ( .A1(n303), .A2(n167), .ZN(n313) );
  CLKBUF_X1 U293 ( .A(n264), .Z(n358) );
  OAI21_X1 U294 ( .B1(n61), .B2(n65), .A(n62), .ZN(n314) );
  OAI21_X1 U295 ( .B1(n310), .B2(n65), .A(n62), .ZN(n2) );
  XNOR2_X1 U296 ( .A(n133), .B(n315), .ZN(n131) );
  XNOR2_X1 U297 ( .A(n138), .B(n135), .ZN(n315) );
  OR2_X1 U298 ( .A1(n121), .A2(n124), .ZN(n316) );
  NOR2_X1 U299 ( .A1(n64), .A2(n310), .ZN(n317) );
  XOR2_X1 U300 ( .A(n167), .B(n184), .Z(n149) );
  BUF_X2 U301 ( .A(n265), .Z(n320) );
  NAND2_X1 U302 ( .A1(n133), .A2(n138), .ZN(n321) );
  NAND2_X1 U303 ( .A1(n133), .A2(n135), .ZN(n322) );
  NAND2_X1 U304 ( .A1(n138), .A2(n135), .ZN(n323) );
  NAND3_X1 U305 ( .A1(n321), .A2(n322), .A3(n323), .ZN(n130) );
  BUF_X1 U306 ( .A(n245), .Z(n360) );
  AND2_X1 U307 ( .A1(n355), .A2(n97), .ZN(product[1]) );
  AOI21_X1 U308 ( .B1(n83), .B2(n308), .A(n339), .ZN(n325) );
  INV_X1 U309 ( .A(n75), .ZN(n326) );
  OAI21_X1 U310 ( .B1(n76), .B2(n325), .A(n77), .ZN(n327) );
  OAI22_X1 U311 ( .A1(n350), .A2(n221), .B1(n220), .B2(n356), .ZN(n328) );
  NAND2_X1 U312 ( .A1(n248), .A2(n256), .ZN(n329) );
  NOR2_X1 U313 ( .A1(n131), .A2(n136), .ZN(n332) );
  NOR2_X1 U314 ( .A1(n131), .A2(n136), .ZN(n69) );
  XOR2_X1 U315 ( .A(n313), .B(n183), .Z(n333) );
  XOR2_X1 U316 ( .A(n145), .B(n333), .Z(n143) );
  NAND2_X1 U317 ( .A1(n145), .A2(n313), .ZN(n334) );
  NAND2_X1 U318 ( .A1(n145), .A2(n183), .ZN(n335) );
  NAND2_X1 U319 ( .A1(n313), .A2(n183), .ZN(n336) );
  NAND3_X1 U320 ( .A1(n334), .A2(n335), .A3(n336), .ZN(n142) );
  CLKBUF_X1 U321 ( .A(n251), .Z(n337) );
  CLKBUF_X1 U322 ( .A(n83), .Z(n338) );
  AND2_X1 U323 ( .A1(n147), .A2(n150), .ZN(n339) );
  INV_X1 U324 ( .A(n158), .ZN(n359) );
  CLKBUF_X1 U325 ( .A(n89), .Z(n341) );
  OAI21_X1 U326 ( .B1(n86), .B2(n84), .A(n85), .ZN(n83) );
  NAND2_X1 U327 ( .A1(n263), .A2(n343), .ZN(n344) );
  NAND2_X1 U328 ( .A1(n342), .A2(a[4]), .ZN(n345) );
  NAND2_X1 U329 ( .A1(n344), .A2(n345), .ZN(n247) );
  INV_X1 U330 ( .A(n263), .ZN(n342) );
  INV_X1 U331 ( .A(a[4]), .ZN(n343) );
  XNOR2_X2 U332 ( .A(n263), .B(a[6]), .ZN(n352) );
  CLKBUF_X1 U333 ( .A(n78), .Z(n346) );
  AOI21_X1 U334 ( .B1(n353), .B2(n83), .A(n339), .ZN(n78) );
  NAND2_X2 U335 ( .A1(n247), .A2(n304), .ZN(n251) );
  NAND2_X1 U336 ( .A1(n246), .A2(n254), .ZN(n348) );
  NAND2_X1 U337 ( .A1(n248), .A2(n256), .ZN(n350) );
  AOI21_X1 U338 ( .B1(n67), .B2(n327), .A(n68), .ZN(n351) );
  AOI21_X1 U339 ( .B1(n67), .B2(n327), .A(n68), .ZN(n1) );
  INV_X1 U340 ( .A(n30), .ZN(n28) );
  NAND2_X1 U341 ( .A1(n103), .A2(n307), .ZN(n9) );
  INV_X1 U342 ( .A(n64), .ZN(n103) );
  INV_X1 U343 ( .A(n18), .ZN(product[15]) );
  INV_X1 U344 ( .A(n31), .ZN(n29) );
  NAND2_X1 U345 ( .A1(n52), .A2(n32), .ZN(n30) );
  NOR2_X1 U346 ( .A1(n332), .A2(n72), .ZN(n67) );
  NAND2_X1 U347 ( .A1(n109), .A2(n341), .ZN(n15) );
  INV_X1 U348 ( .A(n330), .ZN(n109) );
  XNOR2_X1 U349 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U350 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U351 ( .A(n34), .ZN(n99) );
  NAND2_X1 U352 ( .A1(n316), .A2(n62), .ZN(n8) );
  INV_X1 U353 ( .A(n94), .ZN(n92) );
  XNOR2_X1 U354 ( .A(n13), .B(n338), .ZN(product[5]) );
  NAND2_X1 U355 ( .A1(n308), .A2(n82), .ZN(n13) );
  XOR2_X1 U356 ( .A(n86), .B(n14), .Z(product[4]) );
  NAND2_X1 U357 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U358 ( .A(n84), .ZN(n108) );
  NAND2_X1 U359 ( .A1(n105), .A2(n312), .ZN(n11) );
  INV_X1 U360 ( .A(n72), .ZN(n105) );
  XNOR2_X1 U361 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U362 ( .A1(n52), .A2(n51), .ZN(n7) );
  XNOR2_X1 U363 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U364 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U365 ( .A(n41), .ZN(n100) );
  NAND2_X1 U366 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U367 ( .A(n332), .ZN(n104) );
  NAND2_X1 U368 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U369 ( .A(n23), .ZN(n98) );
  AOI21_X1 U370 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U371 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  OAI21_X1 U372 ( .B1(n76), .B2(n78), .A(n77), .ZN(n75) );
  NOR2_X1 U373 ( .A1(n125), .A2(n130), .ZN(n64) );
  NOR2_X1 U374 ( .A1(n41), .A2(n34), .ZN(n32) );
  OAI21_X1 U375 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  INV_X1 U376 ( .A(n50), .ZN(n52) );
  NOR2_X1 U377 ( .A1(n64), .A2(n61), .ZN(n3) );
  NAND2_X1 U378 ( .A1(n125), .A2(n130), .ZN(n65) );
  INV_X1 U379 ( .A(n87), .ZN(n86) );
  OAI21_X1 U380 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U381 ( .A(n51), .ZN(n53) );
  NOR2_X1 U382 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U383 ( .A1(n50), .A2(n41), .ZN(n39) );
  XNOR2_X1 U384 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U385 ( .A1(n354), .A2(n94), .ZN(n16) );
  NAND2_X1 U386 ( .A1(n106), .A2(n77), .ZN(n12) );
  INV_X1 U387 ( .A(n76), .ZN(n106) );
  NOR2_X1 U388 ( .A1(n116), .A2(n115), .ZN(n41) );
  OR2_X1 U389 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U390 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U391 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U392 ( .A(n112), .ZN(n113) );
  NOR2_X1 U393 ( .A1(n117), .A2(n120), .ZN(n50) );
  NOR2_X1 U394 ( .A1(n151), .A2(n152), .ZN(n84) );
  NAND2_X1 U395 ( .A1(n170), .A2(n112), .ZN(n24) );
  XNOR2_X1 U396 ( .A(n187), .B(n175), .ZN(n135) );
  NAND2_X1 U397 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U398 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U399 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U400 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U401 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U402 ( .A1(n151), .A2(n152), .ZN(n85) );
  NAND2_X1 U403 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U404 ( .A1(n143), .A2(n146), .ZN(n77) );
  NAND2_X1 U405 ( .A1(n147), .A2(n150), .ZN(n82) );
  OR2_X1 U406 ( .A1(n200), .A2(n193), .ZN(n354) );
  AND2_X1 U407 ( .A1(n360), .A2(n161), .ZN(n193) );
  OR2_X1 U408 ( .A1(n360), .A2(n260), .ZN(n228) );
  INV_X1 U409 ( .A(n157), .ZN(n178) );
  AND2_X1 U410 ( .A1(n360), .A2(n158), .ZN(n185) );
  INV_X1 U411 ( .A(n118), .ZN(n119) );
  OR2_X1 U412 ( .A1(n360), .A2(n342), .ZN(n219) );
  OR2_X1 U413 ( .A1(n201), .A2(n169), .ZN(n355) );
  INV_X1 U414 ( .A(n163), .ZN(n194) );
  AND2_X1 U415 ( .A1(n360), .A2(n155), .ZN(n177) );
  INV_X1 U416 ( .A(n160), .ZN(n186) );
  INV_X1 U417 ( .A(n154), .ZN(n170) );
  OR2_X1 U418 ( .A1(n360), .A2(n258), .ZN(n210) );
  XNOR2_X1 U419 ( .A(n263), .B(a[6]), .ZN(n254) );
  OR2_X1 U420 ( .A1(n360), .A2(n261), .ZN(n237) );
  NAND2_X1 U421 ( .A1(n246), .A2(n254), .ZN(n250) );
  INV_X1 U422 ( .A(n164), .ZN(n273) );
  AND2_X1 U423 ( .A1(n360), .A2(n164), .ZN(product[0]) );
  AOI21_X1 U424 ( .B1(n354), .B2(n95), .A(n92), .ZN(n90) );
  XNOR2_X1 U425 ( .A(n318), .B(a[2]), .ZN(n256) );
  INV_X1 U426 ( .A(n97), .ZN(n95) );
  XNOR2_X1 U427 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U428 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U429 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U430 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U431 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U432 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U433 ( .A(n262), .B(n360), .ZN(n209) );
  INV_X1 U434 ( .A(n262), .ZN(n258) );
  XNOR2_X1 U435 ( .A(b[1]), .B(n262), .ZN(n208) );
  XOR2_X1 U436 ( .A(a[6]), .B(n262), .Z(n246) );
  OAI22_X1 U437 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  OAI22_X1 U438 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  OAI22_X1 U439 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U440 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U441 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U442 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  OAI22_X1 U443 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OAI22_X1 U444 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  XNOR2_X1 U445 ( .A(n357), .B(a[4]), .ZN(n255) );
  NAND2_X1 U446 ( .A1(n317), .A2(n21), .ZN(n19) );
  NAND2_X1 U447 ( .A1(n317), .A2(n28), .ZN(n26) );
  NAND2_X1 U448 ( .A1(n317), .A2(n39), .ZN(n37) );
  NAND2_X1 U449 ( .A1(n3), .A2(n52), .ZN(n46) );
  INV_X1 U450 ( .A(n3), .ZN(n57) );
  XNOR2_X1 U451 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U452 ( .A1(n200), .A2(n193), .ZN(n94) );
  XNOR2_X1 U453 ( .A(n71), .B(n10), .ZN(product[8]) );
  OAI22_X1 U454 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  NAND2_X1 U455 ( .A1(n131), .A2(n136), .ZN(n70) );
  AOI21_X1 U456 ( .B1(n314), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U457 ( .B1(n314), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U458 ( .B1(n314), .B2(n39), .A(n40), .ZN(n38) );
  INV_X1 U459 ( .A(n314), .ZN(n58) );
  AOI21_X1 U460 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  INV_X1 U461 ( .A(n128), .ZN(n129) );
  OAI21_X1 U462 ( .B1(n326), .B2(n72), .A(n312), .ZN(n71) );
  XOR2_X1 U463 ( .A(n15), .B(n90), .Z(product[3]) );
  OAI21_X1 U464 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NAND2_X1 U465 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI21_X1 U466 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  XNOR2_X1 U467 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U468 ( .A1(n153), .A2(n168), .ZN(n89) );
  NOR2_X1 U469 ( .A1(n153), .A2(n168), .ZN(n88) );
  OAI22_X1 U470 ( .A1(n311), .A2(n217), .B1(n216), .B2(n340), .ZN(n183) );
  OAI22_X1 U471 ( .A1(n337), .A2(n212), .B1(n211), .B2(n340), .ZN(n118) );
  OAI22_X1 U472 ( .A1(n251), .A2(n214), .B1(n213), .B2(n340), .ZN(n180) );
  OAI22_X1 U473 ( .A1(n211), .A2(n337), .B1(n211), .B2(n340), .ZN(n157) );
  OAI22_X1 U474 ( .A1(n251), .A2(n216), .B1(n215), .B2(n340), .ZN(n182) );
  OAI22_X1 U475 ( .A1(n251), .A2(n215), .B1(n214), .B2(n340), .ZN(n181) );
  OAI22_X1 U476 ( .A1(n251), .A2(n213), .B1(n212), .B2(n340), .ZN(n179) );
  INV_X1 U477 ( .A(n255), .ZN(n158) );
  OAI22_X1 U478 ( .A1(n251), .A2(n342), .B1(n219), .B2(n359), .ZN(n167) );
  OAI22_X1 U479 ( .A1(n251), .A2(n218), .B1(n217), .B2(n359), .ZN(n184) );
  XNOR2_X1 U480 ( .A(b[5]), .B(n305), .ZN(n222) );
  XNOR2_X1 U481 ( .A(b[3]), .B(n305), .ZN(n224) );
  XNOR2_X1 U482 ( .A(b[4]), .B(n305), .ZN(n223) );
  XNOR2_X1 U483 ( .A(b[6]), .B(n305), .ZN(n221) );
  XNOR2_X1 U484 ( .A(b[2]), .B(n305), .ZN(n225) );
  INV_X1 U485 ( .A(n305), .ZN(n260) );
  XNOR2_X1 U486 ( .A(b[7]), .B(n305), .ZN(n220) );
  XNOR2_X1 U487 ( .A(n305), .B(n360), .ZN(n227) );
  XNOR2_X1 U488 ( .A(b[1]), .B(n305), .ZN(n226) );
  XOR2_X1 U489 ( .A(n357), .B(a[2]), .Z(n248) );
  OAI22_X1 U490 ( .A1(n202), .A2(n348), .B1(n202), .B2(n352), .ZN(n154) );
  OAI22_X1 U491 ( .A1(n348), .A2(n206), .B1(n205), .B2(n352), .ZN(n173) );
  OAI22_X1 U492 ( .A1(n348), .A2(n203), .B1(n202), .B2(n352), .ZN(n112) );
  OAI22_X1 U493 ( .A1(n348), .A2(n205), .B1(n204), .B2(n352), .ZN(n172) );
  OAI22_X1 U494 ( .A1(n348), .A2(n204), .B1(n203), .B2(n352), .ZN(n171) );
  OAI22_X1 U495 ( .A1(n348), .A2(n208), .B1(n207), .B2(n352), .ZN(n175) );
  OAI22_X1 U496 ( .A1(n348), .A2(n207), .B1(n206), .B2(n352), .ZN(n174) );
  INV_X1 U497 ( .A(n352), .ZN(n155) );
  OAI22_X1 U498 ( .A1(n250), .A2(n258), .B1(n210), .B2(n352), .ZN(n166) );
  OAI22_X1 U499 ( .A1(n250), .A2(n209), .B1(n208), .B2(n352), .ZN(n176) );
  XNOR2_X1 U500 ( .A(b[2]), .B(n331), .ZN(n216) );
  XNOR2_X1 U501 ( .A(b[6]), .B(n347), .ZN(n212) );
  XNOR2_X1 U502 ( .A(b[3]), .B(n331), .ZN(n215) );
  XNOR2_X1 U503 ( .A(b[4]), .B(n331), .ZN(n214) );
  XNOR2_X1 U504 ( .A(b[5]), .B(n347), .ZN(n213) );
  XNOR2_X1 U505 ( .A(b[7]), .B(n347), .ZN(n211) );
  XNOR2_X1 U506 ( .A(n331), .B(n360), .ZN(n218) );
  XNOR2_X1 U507 ( .A(b[1]), .B(n331), .ZN(n217) );
  OAI21_X1 U508 ( .B1(n349), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U509 ( .B1(n349), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U510 ( .B1(n349), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U511 ( .B1(n57), .B2(n1), .A(n58), .ZN(n56) );
  OAI21_X1 U512 ( .B1(n1), .B2(n46), .A(n47), .ZN(n45) );
  XOR2_X1 U513 ( .A(n1), .B(n9), .Z(product[9]) );
  OAI21_X1 U514 ( .B1(n351), .B2(n64), .A(n307), .ZN(n63) );
  XOR2_X1 U515 ( .A(n12), .B(n346), .Z(product[6]) );
  OAI22_X1 U516 ( .A1(n350), .A2(n221), .B1(n220), .B2(n356), .ZN(n128) );
  OAI22_X1 U517 ( .A1(n220), .A2(n329), .B1(n220), .B2(n356), .ZN(n160) );
  OAI22_X1 U518 ( .A1(n350), .A2(n222), .B1(n221), .B2(n356), .ZN(n187) );
  OAI22_X1 U519 ( .A1(n350), .A2(n224), .B1(n223), .B2(n356), .ZN(n189) );
  OAI22_X1 U520 ( .A1(n329), .A2(n225), .B1(n224), .B2(n356), .ZN(n190) );
  OAI22_X1 U521 ( .A1(n329), .A2(n223), .B1(n222), .B2(n356), .ZN(n188) );
  OAI22_X1 U522 ( .A1(n329), .A2(n260), .B1(n228), .B2(n356), .ZN(n168) );
  OAI22_X1 U523 ( .A1(n329), .A2(n226), .B1(n225), .B2(n356), .ZN(n191) );
  XNOR2_X1 U524 ( .A(b[5]), .B(n319), .ZN(n231) );
  XNOR2_X1 U525 ( .A(b[6]), .B(n320), .ZN(n230) );
  XNOR2_X1 U526 ( .A(b[4]), .B(n319), .ZN(n232) );
  INV_X1 U527 ( .A(n356), .ZN(n161) );
  OAI22_X1 U528 ( .A1(n350), .A2(n227), .B1(n226), .B2(n356), .ZN(n192) );
  XNOR2_X1 U529 ( .A(b[7]), .B(n320), .ZN(n229) );
  XNOR2_X1 U530 ( .A(n319), .B(n360), .ZN(n236) );
  XNOR2_X1 U531 ( .A(b[2]), .B(n319), .ZN(n234) );
  XNOR2_X1 U532 ( .A(b[3]), .B(n319), .ZN(n233) );
  INV_X1 U533 ( .A(n320), .ZN(n261) );
  XNOR2_X1 U534 ( .A(b[1]), .B(n319), .ZN(n235) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n103,
         n105, n106, n108, n109, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n163, n164, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n245, n246, n247, n248, n250, n251, n252,
         n253, n254, n255, n256, n258, n259, n260, n261, n262, n263, n264,
         n265, n273, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n357, n358;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n325), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n177), .B(n196), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  BUF_X2 U268 ( .A(n265), .Z(n303) );
  CLKBUF_X1 U269 ( .A(n347), .Z(n304) );
  CLKBUF_X1 U270 ( .A(n263), .Z(n305) );
  CLKBUF_X1 U271 ( .A(n265), .Z(n306) );
  CLKBUF_X1 U272 ( .A(n167), .Z(n307) );
  XNOR2_X1 U273 ( .A(n133), .B(n323), .ZN(n308) );
  NOR2_X1 U274 ( .A1(n121), .A2(n124), .ZN(n309) );
  NAND2_X1 U275 ( .A1(n247), .A2(n255), .ZN(n310) );
  INV_X1 U276 ( .A(n103), .ZN(n311) );
  AND2_X1 U277 ( .A1(n147), .A2(n150), .ZN(n312) );
  INV_X1 U278 ( .A(n82), .ZN(n313) );
  OAI21_X1 U279 ( .B1(n84), .B2(n86), .A(n85), .ZN(n314) );
  CLKBUF_X1 U280 ( .A(n263), .Z(n315) );
  NOR2_X1 U281 ( .A1(n143), .A2(n146), .ZN(n316) );
  NOR2_X1 U282 ( .A1(n143), .A2(n146), .ZN(n76) );
  OAI21_X1 U283 ( .B1(n309), .B2(n65), .A(n62), .ZN(n317) );
  OAI21_X1 U284 ( .B1(n309), .B2(n65), .A(n62), .ZN(n2) );
  CLKBUF_X1 U285 ( .A(n263), .Z(n318) );
  NAND2_X1 U286 ( .A1(n264), .A2(n320), .ZN(n321) );
  NAND2_X1 U287 ( .A1(n319), .A2(a[2]), .ZN(n322) );
  NAND2_X1 U288 ( .A1(n321), .A2(n322), .ZN(n248) );
  INV_X1 U289 ( .A(n264), .ZN(n319) );
  INV_X1 U290 ( .A(a[2]), .ZN(n320) );
  XNOR2_X1 U291 ( .A(n133), .B(n323), .ZN(n131) );
  XNOR2_X1 U292 ( .A(n138), .B(n135), .ZN(n323) );
  OR2_X1 U293 ( .A1(n121), .A2(n124), .ZN(n324) );
  AND2_X1 U294 ( .A1(n184), .A2(n307), .ZN(n325) );
  CLKBUF_X1 U295 ( .A(n263), .Z(n326) );
  NOR2_X1 U296 ( .A1(n339), .A2(n72), .ZN(n67) );
  NAND2_X1 U297 ( .A1(n133), .A2(n138), .ZN(n327) );
  NAND2_X1 U298 ( .A1(n133), .A2(n135), .ZN(n328) );
  NAND2_X1 U299 ( .A1(n138), .A2(n135), .ZN(n329) );
  NAND3_X1 U300 ( .A1(n327), .A2(n328), .A3(n329), .ZN(n130) );
  OR2_X1 U301 ( .A1(n308), .A2(n136), .ZN(n330) );
  XOR2_X1 U302 ( .A(n184), .B(n167), .Z(n149) );
  INV_X1 U303 ( .A(n57), .ZN(n331) );
  CLKBUF_X1 U304 ( .A(n264), .Z(n332) );
  INV_X1 U305 ( .A(n164), .ZN(n273) );
  OR2_X1 U306 ( .A1(n201), .A2(n169), .ZN(n333) );
  XNOR2_X1 U307 ( .A(n352), .B(n334), .ZN(product[9]) );
  AND2_X1 U308 ( .A1(n103), .A2(n65), .ZN(n334) );
  BUF_X1 U309 ( .A(n353), .Z(n335) );
  OR2_X2 U310 ( .A1(n336), .A2(n164), .ZN(n253) );
  XNOR2_X1 U311 ( .A(n265), .B(n164), .ZN(n336) );
  BUF_X2 U312 ( .A(n256), .Z(n357) );
  CLKBUF_X1 U313 ( .A(n303), .Z(n337) );
  NAND2_X1 U314 ( .A1(n255), .A2(n247), .ZN(n338) );
  NAND2_X1 U315 ( .A1(n255), .A2(n247), .ZN(n251) );
  NOR2_X1 U316 ( .A1(n131), .A2(n136), .ZN(n339) );
  NOR2_X1 U317 ( .A1(n308), .A2(n136), .ZN(n69) );
  NAND2_X1 U318 ( .A1(n246), .A2(n254), .ZN(n340) );
  NAND2_X1 U319 ( .A1(n246), .A2(n254), .ZN(n341) );
  NAND2_X1 U320 ( .A1(n246), .A2(n254), .ZN(n250) );
  AOI21_X1 U321 ( .B1(n355), .B2(n314), .A(n313), .ZN(n342) );
  AOI21_X1 U322 ( .B1(n355), .B2(n83), .A(n312), .ZN(n343) );
  AOI21_X1 U323 ( .B1(n355), .B2(n83), .A(n312), .ZN(n78) );
  NAND2_X1 U324 ( .A1(n263), .A2(n344), .ZN(n345) );
  NAND2_X1 U325 ( .A1(n259), .A2(a[4]), .ZN(n346) );
  NAND2_X1 U326 ( .A1(n345), .A2(n346), .ZN(n247) );
  INV_X1 U327 ( .A(a[4]), .ZN(n344) );
  AOI21_X1 U328 ( .B1(n67), .B2(n348), .A(n68), .ZN(n347) );
  AOI21_X1 U329 ( .B1(n67), .B2(n348), .A(n68), .ZN(n352) );
  OAI21_X1 U330 ( .B1(n316), .B2(n342), .A(n77), .ZN(n348) );
  NAND2_X1 U331 ( .A1(n256), .A2(n248), .ZN(n349) );
  XNOR2_X1 U332 ( .A(n264), .B(a[4]), .ZN(n350) );
  XNOR2_X1 U333 ( .A(n264), .B(a[4]), .ZN(n351) );
  AOI21_X1 U334 ( .B1(n67), .B2(n348), .A(n68), .ZN(n1) );
  XNOR2_X1 U335 ( .A(n263), .B(a[6]), .ZN(n353) );
  NOR2_X1 U336 ( .A1(n64), .A2(n61), .ZN(n3) );
  NOR2_X1 U337 ( .A1(n121), .A2(n124), .ZN(n61) );
  BUF_X2 U338 ( .A(n245), .Z(n358) );
  INV_X1 U339 ( .A(n30), .ZN(n28) );
  INV_X1 U340 ( .A(n64), .ZN(n103) );
  INV_X1 U341 ( .A(n18), .ZN(product[15]) );
  AOI21_X1 U342 ( .B1(n317), .B2(n21), .A(n22), .ZN(n20) );
  NAND2_X1 U343 ( .A1(n331), .A2(n21), .ZN(n19) );
  AOI21_X1 U344 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  AOI21_X1 U345 ( .B1(n317), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U346 ( .A(n31), .ZN(n29) );
  NAND2_X1 U347 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U348 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U349 ( .A1(n3), .A2(n39), .ZN(n37) );
  NAND2_X1 U350 ( .A1(n3), .A2(n28), .ZN(n26) );
  INV_X1 U351 ( .A(n317), .ZN(n58) );
  NAND2_X1 U352 ( .A1(n355), .A2(n82), .ZN(n13) );
  NAND2_X1 U353 ( .A1(n324), .A2(n62), .ZN(n8) );
  XNOR2_X1 U354 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U355 ( .A1(n52), .A2(n51), .ZN(n7) );
  INV_X1 U356 ( .A(n3), .ZN(n57) );
  XNOR2_X1 U357 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U358 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U359 ( .A(n41), .ZN(n100) );
  INV_X1 U360 ( .A(n50), .ZN(n52) );
  NAND2_X1 U361 ( .A1(n106), .A2(n77), .ZN(n12) );
  INV_X1 U362 ( .A(n316), .ZN(n106) );
  XNOR2_X1 U363 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U364 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U365 ( .A(n34), .ZN(n99) );
  XNOR2_X1 U366 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U367 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U368 ( .A(n23), .ZN(n98) );
  NAND2_X1 U369 ( .A1(n330), .A2(n70), .ZN(n10) );
  AOI21_X1 U370 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U371 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U372 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U373 ( .A1(n125), .A2(n130), .ZN(n64) );
  XOR2_X1 U374 ( .A(n74), .B(n11), .Z(product[7]) );
  NAND2_X1 U375 ( .A1(n105), .A2(n73), .ZN(n11) );
  INV_X1 U376 ( .A(n72), .ZN(n105) );
  NOR2_X1 U377 ( .A1(n50), .A2(n41), .ZN(n39) );
  NOR2_X1 U378 ( .A1(n41), .A2(n34), .ZN(n32) );
  AOI21_X1 U379 ( .B1(n354), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U380 ( .A(n94), .ZN(n92) );
  OAI21_X1 U381 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U382 ( .A(n51), .ZN(n53) );
  NAND2_X1 U383 ( .A1(n125), .A2(n130), .ZN(n65) );
  AOI21_X1 U384 ( .B1(n317), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U385 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  NAND2_X1 U386 ( .A1(n131), .A2(n136), .ZN(n70) );
  XNOR2_X1 U387 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U388 ( .A1(n354), .A2(n94), .ZN(n16) );
  NOR2_X1 U389 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U390 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U391 ( .A1(n187), .A2(n175), .ZN(n134) );
  XOR2_X1 U392 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U393 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U394 ( .A(n84), .ZN(n108) );
  NOR2_X1 U395 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U396 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U397 ( .A(n112), .ZN(n113) );
  NOR2_X1 U398 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U399 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U400 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U401 ( .A1(n137), .A2(n142), .ZN(n72) );
  INV_X1 U402 ( .A(n97), .ZN(n95) );
  OR2_X1 U403 ( .A1(n200), .A2(n193), .ZN(n354) );
  NAND2_X1 U404 ( .A1(n117), .A2(n120), .ZN(n51) );
  XOR2_X1 U405 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U406 ( .A(n88), .ZN(n109) );
  NAND2_X1 U407 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U408 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U409 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U410 ( .A1(n143), .A2(n146), .ZN(n77) );
  NAND2_X1 U411 ( .A1(n147), .A2(n150), .ZN(n82) );
  OR2_X1 U412 ( .A1(n147), .A2(n150), .ZN(n355) );
  AND2_X1 U413 ( .A1(n358), .A2(n161), .ZN(n193) );
  INV_X1 U414 ( .A(n118), .ZN(n119) );
  AND2_X1 U415 ( .A1(n358), .A2(n158), .ZN(n185) );
  OAI22_X1 U416 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OR2_X1 U417 ( .A1(n358), .A2(n259), .ZN(n219) );
  OAI22_X1 U418 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  AND2_X1 U419 ( .A1(n333), .A2(n97), .ZN(product[1]) );
  INV_X1 U420 ( .A(n163), .ZN(n194) );
  OAI22_X1 U421 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  INV_X1 U422 ( .A(n128), .ZN(n129) );
  AND2_X1 U423 ( .A1(n358), .A2(n155), .ZN(n177) );
  OAI22_X1 U424 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U425 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  NOR2_X1 U426 ( .A1(n151), .A2(n152), .ZN(n84) );
  NOR2_X1 U427 ( .A1(n153), .A2(n168), .ZN(n88) );
  INV_X1 U428 ( .A(n154), .ZN(n170) );
  NAND2_X1 U429 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U430 ( .A1(n358), .A2(n258), .ZN(n210) );
  INV_X1 U431 ( .A(n157), .ZN(n178) );
  XNOR2_X1 U432 ( .A(n263), .B(a[6]), .ZN(n254) );
  XNOR2_X1 U433 ( .A(n264), .B(a[4]), .ZN(n255) );
  OR2_X1 U434 ( .A1(n358), .A2(n260), .ZN(n228) );
  OAI22_X1 U435 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U436 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OAI22_X1 U437 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OR2_X1 U438 ( .A1(n358), .A2(n261), .ZN(n237) );
  XNOR2_X1 U439 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U440 ( .A(b[7]), .B(n262), .ZN(n202) );
  XOR2_X1 U441 ( .A(a[6]), .B(n262), .Z(n246) );
  NAND2_X1 U442 ( .A1(n256), .A2(n248), .ZN(n252) );
  XNOR2_X1 U443 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U444 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U445 ( .A(n262), .B(n358), .ZN(n209) );
  INV_X1 U446 ( .A(n262), .ZN(n258) );
  AND2_X1 U447 ( .A1(n358), .A2(n164), .ZN(product[0]) );
  NAND2_X1 U448 ( .A1(n109), .A2(n89), .ZN(n15) );
  OAI21_X1 U449 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  XNOR2_X1 U450 ( .A(n265), .B(a[2]), .ZN(n256) );
  XOR2_X1 U451 ( .A(n12), .B(n343), .Z(product[6]) );
  XNOR2_X1 U452 ( .A(n303), .B(b[5]), .ZN(n231) );
  XNOR2_X1 U453 ( .A(n303), .B(b[6]), .ZN(n230) );
  XNOR2_X1 U454 ( .A(n337), .B(b[4]), .ZN(n232) );
  XNOR2_X1 U455 ( .A(n337), .B(n358), .ZN(n236) );
  XNOR2_X1 U456 ( .A(n303), .B(b[7]), .ZN(n229) );
  INV_X1 U457 ( .A(n303), .ZN(n261) );
  XNOR2_X1 U458 ( .A(n63), .B(n8), .ZN(product[10]) );
  OAI21_X1 U459 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  INV_X1 U460 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U461 ( .A(n332), .B(b[5]), .ZN(n222) );
  XNOR2_X1 U462 ( .A(n264), .B(b[4]), .ZN(n223) );
  XNOR2_X1 U463 ( .A(n332), .B(b[6]), .ZN(n221) );
  XNOR2_X1 U464 ( .A(n264), .B(b[7]), .ZN(n220) );
  XNOR2_X1 U465 ( .A(n332), .B(n358), .ZN(n227) );
  XNOR2_X1 U466 ( .A(n13), .B(n314), .ZN(product[5]) );
  OAI21_X1 U467 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  NAND2_X1 U468 ( .A1(n200), .A2(n193), .ZN(n94) );
  OAI22_X1 U469 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  INV_X1 U470 ( .A(n160), .ZN(n186) );
  OAI21_X1 U471 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  INV_X1 U472 ( .A(n75), .ZN(n74) );
  XNOR2_X1 U473 ( .A(n264), .B(b[3]), .ZN(n224) );
  XNOR2_X1 U474 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U475 ( .A(n306), .B(b[3]), .ZN(n233) );
  OAI21_X1 U476 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  XNOR2_X1 U477 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U478 ( .A(n332), .B(b[2]), .ZN(n225) );
  XNOR2_X1 U479 ( .A(n306), .B(b[2]), .ZN(n234) );
  NAND2_X1 U480 ( .A1(n201), .A2(n169), .ZN(n97) );
  XNOR2_X1 U481 ( .A(b[1]), .B(n262), .ZN(n208) );
  XNOR2_X1 U482 ( .A(n264), .B(b[1]), .ZN(n226) );
  XNOR2_X1 U483 ( .A(n306), .B(b[1]), .ZN(n235) );
  OAI22_X1 U484 ( .A1(n202), .A2(n340), .B1(n202), .B2(n335), .ZN(n154) );
  OAI22_X1 U485 ( .A1(n341), .A2(n203), .B1(n335), .B2(n202), .ZN(n112) );
  OAI22_X1 U486 ( .A1(n340), .A2(n206), .B1(n335), .B2(n205), .ZN(n173) );
  OAI22_X1 U487 ( .A1(n340), .A2(n205), .B1(n335), .B2(n204), .ZN(n172) );
  OAI22_X1 U488 ( .A1(n341), .A2(n204), .B1(n335), .B2(n203), .ZN(n171) );
  OAI22_X1 U489 ( .A1(n341), .A2(n208), .B1(n353), .B2(n207), .ZN(n175) );
  OAI22_X1 U490 ( .A1(n340), .A2(n207), .B1(n353), .B2(n206), .ZN(n174) );
  INV_X1 U491 ( .A(n353), .ZN(n155) );
  OAI22_X1 U492 ( .A1(n250), .A2(n258), .B1(n210), .B2(n353), .ZN(n166) );
  OAI22_X1 U493 ( .A1(n250), .A2(n209), .B1(n353), .B2(n208), .ZN(n176) );
  XNOR2_X1 U494 ( .A(n315), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U495 ( .A(n305), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U496 ( .A(n326), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U497 ( .A(n326), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U498 ( .A(n318), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U499 ( .A(n305), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U500 ( .A(n305), .B(n358), .ZN(n218) );
  INV_X1 U501 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U502 ( .A(n263), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U503 ( .A(n71), .B(n10), .ZN(product[8]) );
  INV_X1 U504 ( .A(n87), .ZN(n86) );
  OAI21_X1 U505 ( .B1(n352), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U506 ( .B1(n352), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U507 ( .B1(n304), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U508 ( .B1(n347), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U509 ( .B1(n347), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U510 ( .B1(n1), .B2(n311), .A(n65), .ZN(n63) );
  OAI22_X1 U511 ( .A1(n310), .A2(n217), .B1(n216), .B2(n350), .ZN(n183) );
  OAI22_X1 U512 ( .A1(n338), .A2(n212), .B1(n211), .B2(n351), .ZN(n118) );
  OAI22_X1 U513 ( .A1(n211), .A2(n310), .B1(n211), .B2(n350), .ZN(n157) );
  OAI22_X1 U514 ( .A1(n310), .A2(n213), .B1(n212), .B2(n351), .ZN(n179) );
  OAI22_X1 U515 ( .A1(n338), .A2(n214), .B1(n213), .B2(n350), .ZN(n180) );
  OAI22_X1 U516 ( .A1(n310), .A2(n216), .B1(n215), .B2(n351), .ZN(n182) );
  OAI22_X1 U517 ( .A1(n338), .A2(n215), .B1(n214), .B2(n350), .ZN(n181) );
  INV_X1 U518 ( .A(n351), .ZN(n158) );
  OAI22_X1 U519 ( .A1(n251), .A2(n259), .B1(n219), .B2(n350), .ZN(n167) );
  OAI22_X1 U520 ( .A1(n251), .A2(n218), .B1(n217), .B2(n351), .ZN(n184) );
  NAND2_X1 U521 ( .A1(n153), .A2(n168), .ZN(n89) );
  OAI22_X1 U522 ( .A1(n349), .A2(n221), .B1(n220), .B2(n357), .ZN(n128) );
  OAI22_X1 U523 ( .A1(n252), .A2(n222), .B1(n221), .B2(n357), .ZN(n187) );
  OAI22_X1 U524 ( .A1(n349), .A2(n224), .B1(n223), .B2(n357), .ZN(n189) );
  OAI22_X1 U525 ( .A1(n252), .A2(n225), .B1(n224), .B2(n357), .ZN(n190) );
  OAI22_X1 U526 ( .A1(n252), .A2(n223), .B1(n222), .B2(n357), .ZN(n188) );
  OAI22_X1 U527 ( .A1(n220), .A2(n349), .B1(n220), .B2(n357), .ZN(n160) );
  OAI22_X1 U528 ( .A1(n252), .A2(n260), .B1(n228), .B2(n357), .ZN(n168) );
  OAI22_X1 U529 ( .A1(n252), .A2(n226), .B1(n225), .B2(n357), .ZN(n191) );
  OAI22_X1 U530 ( .A1(n349), .A2(n227), .B1(n226), .B2(n357), .ZN(n192) );
  INV_X1 U531 ( .A(n357), .ZN(n161) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_3_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n21, n22, n26, n27, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n51, n52, n54, n56,
         n57, n58, n60, n62, n63, n64, n65, n66, n68, n70, n71, n72, n73, n74,
         n76, n78, n79, n80, n81, n82, n84, n86, n87, n89, n92, n95, n99, n101,
         n103, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193;

  OR2_X2 U125 ( .A1(A[9]), .A2(B[9]), .ZN(n192) );
  CLKBUF_X1 U126 ( .A(n183), .Z(n160) );
  CLKBUF_X1 U127 ( .A(B[12]), .Z(n161) );
  OR2_X1 U128 ( .A1(A[14]), .A2(B[14]), .ZN(n186) );
  AND2_X1 U129 ( .A1(B[14]), .A2(A[14]), .ZN(n163) );
  AND2_X1 U130 ( .A1(B[9]), .A2(A[9]), .ZN(n162) );
  INV_X4 U131 ( .A(n162), .ZN(n51) );
  INV_X4 U132 ( .A(n163), .ZN(n26) );
  CLKBUF_X1 U133 ( .A(A[12]), .Z(n164) );
  NOR2_X2 U134 ( .A1(B[10]), .A2(A[10]), .ZN(n42) );
  OAI21_X1 U135 ( .B1(n74), .B2(n72), .A(n73), .ZN(n165) );
  CLKBUF_X1 U136 ( .A(n56), .Z(n170) );
  XNOR2_X1 U137 ( .A(n44), .B(n166), .ZN(SUM[10]) );
  AND2_X1 U138 ( .A1(n95), .A2(n43), .ZN(n166) );
  AOI21_X1 U139 ( .B1(n190), .B2(n79), .A(n76), .ZN(n167) );
  BUF_X1 U140 ( .A(n181), .Z(n168) );
  CLKBUF_X1 U141 ( .A(n43), .Z(n169) );
  BUF_X1 U142 ( .A(n40), .Z(n171) );
  CLKBUF_X1 U143 ( .A(B[11]), .Z(n172) );
  BUF_X1 U144 ( .A(n33), .Z(n173) );
  CLKBUF_X1 U145 ( .A(A[11]), .Z(n174) );
  NAND2_X1 U146 ( .A1(B[10]), .A2(A[10]), .ZN(n43) );
  OR2_X1 U147 ( .A1(B[0]), .A2(A[0]), .ZN(n175) );
  AND2_X1 U148 ( .A1(n175), .A2(n89), .ZN(SUM[0]) );
  BUF_X1 U149 ( .A(n35), .Z(n177) );
  OR2_X1 U150 ( .A1(n183), .A2(n35), .ZN(n178) );
  AOI21_X1 U151 ( .B1(n45), .B2(n37), .A(n38), .ZN(n179) );
  AOI21_X1 U152 ( .B1(n45), .B2(n37), .A(n38), .ZN(n1) );
  OR2_X1 U153 ( .A1(n161), .A2(n164), .ZN(n180) );
  CLKBUF_X1 U154 ( .A(n36), .Z(n181) );
  NOR2_X1 U155 ( .A1(A[12]), .A2(B[12]), .ZN(n35) );
  NOR2_X1 U156 ( .A1(B[11]), .A2(A[11]), .ZN(n182) );
  NOR2_X1 U157 ( .A1(B[13]), .A2(A[13]), .ZN(n183) );
  INV_X1 U158 ( .A(n62), .ZN(n60) );
  INV_X1 U159 ( .A(n42), .ZN(n95) );
  NAND2_X1 U160 ( .A1(n92), .A2(n173), .ZN(n4) );
  INV_X1 U161 ( .A(n160), .ZN(n92) );
  XNOR2_X1 U162 ( .A(n184), .B(n52), .ZN(SUM[9]) );
  AND2_X1 U163 ( .A1(n192), .A2(n51), .ZN(n184) );
  XNOR2_X1 U164 ( .A(n165), .B(n12), .ZN(SUM[5]) );
  NAND2_X1 U165 ( .A1(n99), .A2(n65), .ZN(n11) );
  INV_X1 U166 ( .A(n64), .ZN(n99) );
  NAND2_X1 U167 ( .A1(n180), .A2(n181), .ZN(n5) );
  NAND2_X1 U168 ( .A1(n187), .A2(n62), .ZN(n10) );
  INV_X1 U169 ( .A(n78), .ZN(n76) );
  NOR2_X1 U170 ( .A1(A[13]), .A2(B[13]), .ZN(n32) );
  NAND2_X1 U171 ( .A1(n185), .A2(n19), .ZN(n2) );
  NAND2_X1 U172 ( .A1(B[6]), .A2(A[6]), .ZN(n65) );
  OR2_X1 U173 ( .A1(B[15]), .A2(A[15]), .ZN(n185) );
  NOR2_X1 U174 ( .A1(B[6]), .A2(A[6]), .ZN(n64) );
  XNOR2_X1 U175 ( .A(n41), .B(n6), .ZN(SUM[11]) );
  NAND2_X1 U176 ( .A1(n193), .A2(n171), .ZN(n6) );
  OR2_X1 U177 ( .A1(B[7]), .A2(A[7]), .ZN(n187) );
  OR2_X1 U178 ( .A1(B[5]), .A2(A[5]), .ZN(n188) );
  OR2_X1 U179 ( .A1(B[8]), .A2(A[8]), .ZN(n189) );
  XNOR2_X1 U180 ( .A(n14), .B(n79), .ZN(SUM[3]) );
  NAND2_X1 U181 ( .A1(n190), .A2(n78), .ZN(n14) );
  NAND2_X1 U182 ( .A1(n101), .A2(n73), .ZN(n13) );
  INV_X1 U183 ( .A(n72), .ZN(n101) );
  OAI21_X1 U184 ( .B1(n82), .B2(n80), .A(n81), .ZN(n79) );
  XOR2_X1 U185 ( .A(n15), .B(n82), .Z(SUM[2]) );
  NAND2_X1 U186 ( .A1(n103), .A2(n81), .ZN(n15) );
  INV_X1 U187 ( .A(n80), .ZN(n103) );
  NOR2_X1 U188 ( .A1(B[4]), .A2(A[4]), .ZN(n72) );
  NAND2_X1 U189 ( .A1(B[4]), .A2(A[4]), .ZN(n73) );
  OR2_X1 U190 ( .A1(B[3]), .A2(A[3]), .ZN(n190) );
  AOI21_X1 U191 ( .B1(n191), .B2(n87), .A(n84), .ZN(n82) );
  INV_X1 U192 ( .A(n86), .ZN(n84) );
  NOR2_X1 U193 ( .A1(B[2]), .A2(A[2]), .ZN(n80) );
  NAND2_X1 U194 ( .A1(B[2]), .A2(A[2]), .ZN(n81) );
  XNOR2_X1 U195 ( .A(n16), .B(n87), .ZN(SUM[1]) );
  NAND2_X1 U196 ( .A1(n191), .A2(n86), .ZN(n16) );
  OR2_X1 U197 ( .A1(B[1]), .A2(A[1]), .ZN(n191) );
  INV_X1 U198 ( .A(n89), .ZN(n87) );
  NAND2_X1 U199 ( .A1(B[1]), .A2(A[1]), .ZN(n86) );
  NAND2_X1 U200 ( .A1(B[0]), .A2(A[0]), .ZN(n89) );
  XNOR2_X1 U201 ( .A(n9), .B(n57), .ZN(SUM[8]) );
  INV_X1 U202 ( .A(n70), .ZN(n68) );
  NAND2_X1 U203 ( .A1(n188), .A2(n70), .ZN(n12) );
  NAND2_X1 U204 ( .A1(B[5]), .A2(A[5]), .ZN(n70) );
  AOI21_X1 U205 ( .B1(n190), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U206 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  OAI21_X1 U207 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  AOI21_X1 U208 ( .B1(n71), .B2(n188), .A(n68), .ZN(n66) );
  NAND2_X1 U209 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NAND2_X1 U210 ( .A1(n186), .A2(n26), .ZN(n3) );
  INV_X1 U211 ( .A(n58), .ZN(n57) );
  AOI21_X1 U212 ( .B1(n63), .B2(n187), .A(n60), .ZN(n58) );
  OR2_X1 U213 ( .A1(n172), .A2(n174), .ZN(n193) );
  XNOR2_X1 U214 ( .A(n63), .B(n10), .ZN(SUM[7]) );
  OAI21_X1 U215 ( .B1(n64), .B2(n66), .A(n65), .ZN(n63) );
  NOR2_X1 U216 ( .A1(n183), .A2(n35), .ZN(n30) );
  AOI21_X1 U217 ( .B1(n189), .B2(n57), .A(n54), .ZN(n52) );
  NAND2_X1 U218 ( .A1(n189), .A2(n170), .ZN(n9) );
  NAND2_X1 U219 ( .A1(B[8]), .A2(A[8]), .ZN(n56) );
  INV_X1 U220 ( .A(n56), .ZN(n54) );
  INV_X1 U221 ( .A(n31), .ZN(n29) );
  NAND2_X1 U222 ( .A1(A[13]), .A2(B[13]), .ZN(n33) );
  NAND2_X1 U223 ( .A1(B[11]), .A2(A[11]), .ZN(n40) );
  NOR2_X1 U224 ( .A1(B[11]), .A2(A[11]), .ZN(n39) );
  XOR2_X1 U225 ( .A(n167), .B(n13), .Z(SUM[4]) );
  XOR2_X1 U226 ( .A(n11), .B(n66), .Z(SUM[6]) );
  NAND2_X1 U227 ( .A1(B[3]), .A2(A[3]), .ZN(n78) );
  NAND2_X1 U228 ( .A1(n192), .A2(n189), .ZN(n46) );
  AOI21_X1 U229 ( .B1(n192), .B2(n54), .A(n162), .ZN(n47) );
  OAI21_X1 U230 ( .B1(n39), .B2(n43), .A(n40), .ZN(n38) );
  OAI21_X1 U231 ( .B1(n44), .B2(n42), .A(n169), .ZN(n41) );
  INV_X1 U232 ( .A(n45), .ZN(n44) );
  XNOR2_X1 U233 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  OAI21_X1 U234 ( .B1(n46), .B2(n58), .A(n47), .ZN(n45) );
  NOR2_X1 U235 ( .A1(n182), .A2(n42), .ZN(n37) );
  XNOR2_X1 U236 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U237 ( .A1(n30), .A2(n186), .ZN(n21) );
  AOI21_X1 U238 ( .B1(n31), .B2(n186), .A(n163), .ZN(n22) );
  OAI21_X1 U239 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U240 ( .A1(A[12]), .A2(B[12]), .ZN(n36) );
  XNOR2_X1 U241 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XOR2_X1 U242 ( .A(n179), .B(n5), .Z(SUM[12]) );
  OAI21_X1 U243 ( .B1(n179), .B2(n178), .A(n29), .ZN(n27) );
  OAI21_X1 U244 ( .B1(n1), .B2(n177), .A(n168), .ZN(n34) );
  OAI21_X1 U245 ( .B1(n1), .B2(n21), .A(n22), .ZN(n20) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_3 ( .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;


  recursive_add_layer_INPUT_SCALE2_WIDTH16_3_DW01_add_2 add_56 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM(out) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_3_DW01_add_4 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34,
         n35, n36, n37, n38, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n59, n60, n62, n64, n65, n66, n68, n70, n71,
         n72, n73, n74, n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89,
         n91, n93, n96, n97, n98, n102, n104, n106, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186;

  BUF_X1 U127 ( .A(n43), .Z(n162) );
  CLKBUF_X1 U128 ( .A(n37), .Z(n166) );
  NOR2_X1 U129 ( .A1(B[12]), .A2(A[12]), .ZN(n163) );
  BUF_X1 U130 ( .A(n74), .Z(n164) );
  INV_X1 U131 ( .A(n168), .ZN(n59) );
  AND2_X1 U132 ( .A1(B[8]), .A2(A[8]), .ZN(n168) );
  CLKBUF_X1 U133 ( .A(n184), .Z(n165) );
  INV_X1 U134 ( .A(n36), .ZN(n167) );
  OR2_X2 U135 ( .A1(B[8]), .A2(A[8]), .ZN(n184) );
  OR2_X1 U136 ( .A1(B[12]), .A2(A[12]), .ZN(n169) );
  AOI21_X1 U137 ( .B1(n184), .B2(n62), .A(n168), .ZN(n170) );
  OR2_X1 U138 ( .A1(A[13]), .A2(B[13]), .ZN(n171) );
  AND2_X1 U139 ( .A1(n180), .A2(n91), .ZN(SUM[0]) );
  XNOR2_X1 U140 ( .A(n53), .B(n173), .ZN(SUM[9]) );
  NAND2_X1 U141 ( .A1(n98), .A2(n51), .ZN(n173) );
  AOI21_X1 U142 ( .B1(n185), .B2(n71), .A(n68), .ZN(n174) );
  CLKBUF_X1 U143 ( .A(n1), .Z(n175) );
  NOR2_X1 U144 ( .A1(B[10]), .A2(A[10]), .ZN(n176) );
  NOR2_X1 U145 ( .A1(A[10]), .A2(B[10]), .ZN(n47) );
  AOI21_X1 U146 ( .B1(n178), .B2(n45), .A(n46), .ZN(n179) );
  NOR2_X1 U147 ( .A1(A[9]), .A2(B[9]), .ZN(n50) );
  XNOR2_X1 U148 ( .A(n1), .B(n177), .ZN(SUM[11]) );
  AND2_X1 U149 ( .A1(n96), .A2(n162), .ZN(n177) );
  INV_X1 U150 ( .A(n50), .ZN(n98) );
  OAI21_X1 U151 ( .B1(n54), .B2(n174), .A(n55), .ZN(n178) );
  AOI21_X1 U152 ( .B1(n178), .B2(n45), .A(n46), .ZN(n1) );
  OR2_X1 U153 ( .A1(B[7]), .A2(A[7]), .ZN(n182) );
  OR2_X1 U154 ( .A1(B[0]), .A2(A[0]), .ZN(n180) );
  INV_X1 U155 ( .A(n38), .ZN(n36) );
  NAND2_X1 U156 ( .A1(n102), .A2(n73), .ZN(n12) );
  OAI21_X1 U157 ( .B1(n163), .B2(n43), .A(n40), .ZN(n38) );
  INV_X1 U158 ( .A(n42), .ZN(n96) );
  NAND2_X1 U159 ( .A1(n169), .A2(n40), .ZN(n5) );
  NAND2_X1 U160 ( .A1(n171), .A2(n33), .ZN(n4) );
  INV_X1 U161 ( .A(n70), .ZN(n68) );
  XNOR2_X1 U162 ( .A(n49), .B(n7), .ZN(SUM[10]) );
  NAND2_X1 U163 ( .A1(n97), .A2(n48), .ZN(n7) );
  INV_X1 U164 ( .A(n176), .ZN(n97) );
  XNOR2_X1 U165 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U166 ( .A1(n93), .A2(n26), .ZN(n3) );
  NOR2_X1 U167 ( .A1(n32), .A2(n25), .ZN(n23) );
  XOR2_X1 U168 ( .A(n60), .B(n9), .Z(SUM[8]) );
  AOI21_X1 U169 ( .B1(n65), .B2(n182), .A(n62), .ZN(n60) );
  INV_X1 U170 ( .A(n33), .ZN(n31) );
  NAND2_X1 U171 ( .A1(n181), .A2(n19), .ZN(n2) );
  NAND2_X1 U172 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NOR2_X1 U173 ( .A1(n42), .A2(n163), .ZN(n37) );
  XNOR2_X1 U174 ( .A(n10), .B(n65), .ZN(SUM[7]) );
  NAND2_X1 U175 ( .A1(n182), .A2(n64), .ZN(n10) );
  OAI21_X1 U176 ( .B1(n47), .B2(n51), .A(n48), .ZN(n46) );
  AOI21_X1 U177 ( .B1(n167), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U178 ( .A(n64), .ZN(n62) );
  OR2_X1 U179 ( .A1(B[15]), .A2(A[15]), .ZN(n181) );
  NAND2_X1 U180 ( .A1(n185), .A2(n70), .ZN(n11) );
  XNOR2_X1 U181 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  NAND2_X1 U182 ( .A1(n186), .A2(n78), .ZN(n13) );
  OAI21_X1 U183 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  XOR2_X1 U184 ( .A(n14), .B(n82), .Z(SUM[3]) );
  NAND2_X1 U185 ( .A1(n104), .A2(n81), .ZN(n14) );
  INV_X1 U186 ( .A(n80), .ZN(n104) );
  NAND2_X1 U187 ( .A1(A[11]), .A2(B[11]), .ZN(n43) );
  AOI21_X1 U188 ( .B1(n186), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U189 ( .A(n78), .ZN(n76) );
  NOR2_X1 U190 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  NOR2_X1 U191 ( .A1(A[11]), .A2(B[11]), .ZN(n42) );
  OR2_X1 U192 ( .A1(B[2]), .A2(A[2]), .ZN(n183) );
  NAND2_X1 U193 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  NOR2_X1 U194 ( .A1(A[13]), .A2(B[13]), .ZN(n32) );
  NAND2_X1 U195 ( .A1(A[13]), .A2(B[13]), .ZN(n33) );
  NAND2_X1 U196 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U197 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  OR2_X1 U198 ( .A1(B[6]), .A2(A[6]), .ZN(n185) );
  XNOR2_X1 U199 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U200 ( .A1(n183), .A2(n86), .ZN(n15) );
  NOR2_X1 U201 ( .A1(A[3]), .A2(B[3]), .ZN(n80) );
  AOI21_X1 U202 ( .B1(n87), .B2(n183), .A(n84), .ZN(n82) );
  INV_X1 U203 ( .A(n86), .ZN(n84) );
  NAND2_X1 U204 ( .A1(A[3]), .A2(B[3]), .ZN(n81) );
  OR2_X1 U205 ( .A1(B[4]), .A2(A[4]), .ZN(n186) );
  NAND2_X1 U206 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  XOR2_X1 U207 ( .A(n16), .B(n91), .Z(SUM[1]) );
  NAND2_X1 U208 ( .A1(n106), .A2(n89), .ZN(n16) );
  INV_X1 U209 ( .A(n88), .ZN(n106) );
  OAI21_X1 U210 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U211 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U212 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  NAND2_X1 U213 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  NOR2_X1 U214 ( .A1(n176), .A2(n50), .ZN(n45) );
  NAND2_X1 U215 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  NAND2_X1 U216 ( .A1(n23), .A2(n166), .ZN(n21) );
  INV_X1 U217 ( .A(n37), .ZN(n35) );
  OAI21_X1 U218 ( .B1(n54), .B2(n174), .A(n170), .ZN(n53) );
  INV_X1 U219 ( .A(n66), .ZN(n65) );
  NAND2_X1 U220 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  NAND2_X1 U221 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  NOR2_X1 U222 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  INV_X1 U223 ( .A(n25), .ZN(n93) );
  OAI21_X1 U224 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  XNOR2_X1 U225 ( .A(n11), .B(n71), .ZN(SUM[6]) );
  AOI21_X1 U226 ( .B1(n185), .B2(n71), .A(n68), .ZN(n66) );
  OAI21_X1 U227 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  XNOR2_X1 U228 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U229 ( .A1(A[7]), .A2(B[7]), .ZN(n64) );
  NAND2_X1 U230 ( .A1(n37), .A2(n171), .ZN(n28) );
  AOI21_X1 U231 ( .B1(n38), .B2(n171), .A(n31), .ZN(n29) );
  INV_X1 U232 ( .A(n72), .ZN(n102) );
  XNOR2_X1 U233 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U234 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  XNOR2_X1 U235 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  XOR2_X1 U236 ( .A(n12), .B(n164), .Z(SUM[5]) );
  INV_X1 U237 ( .A(n53), .ZN(n52) );
  OAI21_X1 U238 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X1 U239 ( .B1(n175), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U240 ( .B1(n1), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U241 ( .B1(n179), .B2(n35), .A(n36), .ZN(n34) );
  OAI21_X1 U242 ( .B1(n42), .B2(n179), .A(n162), .ZN(n41) );
  NAND2_X1 U243 ( .A1(n165), .A2(n59), .ZN(n9) );
  AOI21_X1 U244 ( .B1(n184), .B2(n62), .A(n168), .ZN(n55) );
  NAND2_X1 U245 ( .A1(n184), .A2(n182), .ZN(n54) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_3_DW01_add_5 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n59, n60, n64, n65, n66, n68, n70, n71, n72,
         n73, n74, n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89, n91,
         n93, n94, n96, n97, n102, n104, n106, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188;

  CLKBUF_X1 U127 ( .A(B[12]), .Z(n162) );
  AOI21_X1 U128 ( .B1(n188), .B2(n175), .A(n165), .ZN(n163) );
  OAI21_X1 U129 ( .B1(n54), .B2(n66), .A(n163), .ZN(n164) );
  AND2_X1 U130 ( .A1(B[8]), .A2(A[8]), .ZN(n165) );
  INV_X4 U131 ( .A(n165), .ZN(n59) );
  CLKBUF_X1 U132 ( .A(n48), .Z(n166) );
  NOR2_X1 U133 ( .A1(B[11]), .A2(A[11]), .ZN(n167) );
  NOR2_X1 U134 ( .A1(B[11]), .A2(A[11]), .ZN(n42) );
  NOR2_X1 U135 ( .A1(n179), .A2(n50), .ZN(n168) );
  CLKBUF_X1 U136 ( .A(n51), .Z(n169) );
  OR2_X1 U137 ( .A1(n167), .A2(n39), .ZN(n170) );
  NOR2_X1 U138 ( .A1(B[12]), .A2(A[12]), .ZN(n171) );
  INV_X1 U139 ( .A(n36), .ZN(n172) );
  AND2_X1 U140 ( .A1(B[7]), .A2(A[7]), .ZN(n175) );
  INV_X1 U141 ( .A(n175), .ZN(n64) );
  AND2_X1 U142 ( .A1(n182), .A2(n91), .ZN(SUM[0]) );
  OR2_X1 U143 ( .A1(B[9]), .A2(A[9]), .ZN(n174) );
  OAI21_X1 U144 ( .B1(n54), .B2(n66), .A(n55), .ZN(n53) );
  XNOR2_X1 U145 ( .A(n164), .B(n181), .ZN(SUM[9]) );
  OR2_X1 U146 ( .A1(A[12]), .A2(n162), .ZN(n176) );
  XNOR2_X1 U147 ( .A(n1), .B(n177), .ZN(SUM[11]) );
  AND2_X1 U148 ( .A1(n96), .A2(n43), .ZN(n177) );
  CLKBUF_X1 U149 ( .A(n180), .Z(n178) );
  NOR2_X1 U150 ( .A1(B[10]), .A2(A[10]), .ZN(n179) );
  NOR2_X1 U151 ( .A1(B[10]), .A2(A[10]), .ZN(n47) );
  AOI21_X1 U152 ( .B1(n45), .B2(n53), .A(n46), .ZN(n180) );
  AOI21_X1 U153 ( .B1(n168), .B2(n53), .A(n46), .ZN(n1) );
  NAND2_X1 U154 ( .A1(n174), .A2(n51), .ZN(n181) );
  OR2_X1 U155 ( .A1(B[0]), .A2(A[0]), .ZN(n182) );
  NAND2_X1 U156 ( .A1(n102), .A2(n73), .ZN(n12) );
  INV_X1 U157 ( .A(n72), .ZN(n102) );
  XNOR2_X1 U158 ( .A(n11), .B(n71), .ZN(SUM[6]) );
  NAND2_X1 U159 ( .A1(n186), .A2(n70), .ZN(n11) );
  INV_X1 U160 ( .A(n70), .ZN(n68) );
  NAND2_X1 U161 ( .A1(n94), .A2(n33), .ZN(n4) );
  NAND2_X1 U162 ( .A1(n183), .A2(n19), .ZN(n2) );
  NAND2_X1 U163 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  OAI21_X1 U164 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  XNOR2_X1 U165 ( .A(n49), .B(n7), .ZN(SUM[10]) );
  NAND2_X1 U166 ( .A1(n176), .A2(n40), .ZN(n5) );
  NAND2_X1 U167 ( .A1(n93), .A2(n26), .ZN(n3) );
  XNOR2_X1 U168 ( .A(n10), .B(n65), .ZN(SUM[7]) );
  AOI21_X1 U169 ( .B1(n65), .B2(n185), .A(n175), .ZN(n60) );
  OR2_X1 U170 ( .A1(B[15]), .A2(A[15]), .ZN(n183) );
  INV_X1 U171 ( .A(n33), .ZN(n31) );
  AOI21_X1 U172 ( .B1(n187), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U173 ( .A(n78), .ZN(n76) );
  XOR2_X1 U174 ( .A(n14), .B(n82), .Z(SUM[3]) );
  NAND2_X1 U175 ( .A1(n104), .A2(n81), .ZN(n14) );
  INV_X1 U176 ( .A(n80), .ZN(n104) );
  NOR2_X1 U177 ( .A1(A[12]), .A2(B[12]), .ZN(n39) );
  NOR2_X1 U178 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  OAI21_X1 U179 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  OR2_X1 U180 ( .A1(B[2]), .A2(A[2]), .ZN(n184) );
  NAND2_X1 U181 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  OR2_X1 U182 ( .A1(A[7]), .A2(B[7]), .ZN(n185) );
  NAND2_X1 U183 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U184 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  OR2_X1 U185 ( .A1(B[6]), .A2(A[6]), .ZN(n186) );
  XNOR2_X1 U186 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  NAND2_X1 U187 ( .A1(n187), .A2(n78), .ZN(n13) );
  AOI21_X1 U188 ( .B1(n87), .B2(n184), .A(n84), .ZN(n82) );
  INV_X1 U189 ( .A(n86), .ZN(n84) );
  NAND2_X1 U190 ( .A1(B[3]), .A2(A[3]), .ZN(n81) );
  NOR2_X1 U191 ( .A1(B[3]), .A2(A[3]), .ZN(n80) );
  NAND2_X1 U192 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  OR2_X1 U193 ( .A1(B[4]), .A2(A[4]), .ZN(n187) );
  XNOR2_X1 U194 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U195 ( .A1(n184), .A2(n86), .ZN(n15) );
  OAI21_X1 U196 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U197 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U198 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  XOR2_X1 U199 ( .A(n16), .B(n91), .Z(SUM[1]) );
  NAND2_X1 U200 ( .A1(n106), .A2(n89), .ZN(n16) );
  INV_X1 U201 ( .A(n88), .ZN(n106) );
  NAND2_X1 U202 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  NAND2_X1 U203 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  NOR2_X1 U204 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  NOR2_X1 U205 ( .A1(n167), .A2(n39), .ZN(n37) );
  INV_X1 U206 ( .A(n42), .ZN(n96) );
  NAND2_X1 U207 ( .A1(n97), .A2(n166), .ZN(n7) );
  OR2_X1 U208 ( .A1(B[8]), .A2(A[8]), .ZN(n188) );
  NOR2_X1 U209 ( .A1(n32), .A2(n25), .ZN(n23) );
  INV_X1 U210 ( .A(n32), .ZN(n94) );
  NOR2_X1 U211 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND2_X1 U212 ( .A1(n37), .A2(n23), .ZN(n21) );
  NOR2_X1 U213 ( .A1(B[9]), .A2(A[9]), .ZN(n50) );
  NAND2_X1 U214 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  NAND2_X1 U215 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  NAND2_X1 U216 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  AOI21_X1 U217 ( .B1(n186), .B2(n71), .A(n68), .ZN(n66) );
  INV_X1 U218 ( .A(n66), .ZN(n65) );
  XOR2_X1 U219 ( .A(n12), .B(n74), .Z(SUM[5]) );
  XOR2_X1 U220 ( .A(n60), .B(n9), .Z(SUM[8]) );
  OAI21_X1 U221 ( .B1(n52), .B2(n50), .A(n169), .ZN(n49) );
  NAND2_X1 U222 ( .A1(n185), .A2(n64), .ZN(n10) );
  OAI21_X1 U223 ( .B1(n43), .B2(n171), .A(n40), .ZN(n38) );
  AOI21_X1 U224 ( .B1(n23), .B2(n172), .A(n24), .ZN(n22) );
  INV_X1 U225 ( .A(n38), .ZN(n36) );
  XNOR2_X1 U226 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  INV_X1 U227 ( .A(n25), .ZN(n93) );
  OAI21_X1 U228 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  XNOR2_X1 U229 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  NAND2_X1 U230 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  XNOR2_X1 U231 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U232 ( .A1(n37), .A2(n94), .ZN(n28) );
  AOI21_X1 U233 ( .B1(n38), .B2(n94), .A(n31), .ZN(n29) );
  NAND2_X1 U234 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  XNOR2_X1 U235 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  INV_X1 U236 ( .A(n179), .ZN(n97) );
  NOR2_X1 U237 ( .A1(n179), .A2(n50), .ZN(n45) );
  OAI21_X1 U238 ( .B1(n47), .B2(n51), .A(n48), .ZN(n46) );
  INV_X1 U239 ( .A(n164), .ZN(n52) );
  OAI21_X1 U240 ( .B1(n178), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U241 ( .B1(n180), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U242 ( .B1(n1), .B2(n170), .A(n36), .ZN(n34) );
  OAI21_X1 U243 ( .B1(n180), .B2(n167), .A(n43), .ZN(n41) );
  NAND2_X1 U244 ( .A1(n188), .A2(n59), .ZN(n9) );
  AOI21_X1 U245 ( .B1(n188), .B2(n175), .A(n165), .ZN(n55) );
  NAND2_X1 U246 ( .A1(n188), .A2(n185), .ZN(n54) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_3 ( .in({\in[3][15] , 
        \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , \in[3][10] , 
        \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , \in[3][5] , \in[3][4] , 
        \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , \in[2][15] , 
        \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , \in[2][10] , 
        \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , \in[2][5] , \in[2][4] , 
        \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , \in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \genblk1.inter[1][15] , \genblk1.inter[1][14] ,
         \genblk1.inter[1][13] , \genblk1.inter[1][12] ,
         \genblk1.inter[1][11] , \genblk1.inter[1][10] , \genblk1.inter[1][9] ,
         \genblk1.inter[1][8] , \genblk1.inter[1][7] , \genblk1.inter[1][6] ,
         \genblk1.inter[1][5] , \genblk1.inter[1][4] , \genblk1.inter[1][3] ,
         \genblk1.inter[1][2] , \genblk1.inter[1][1] , \genblk1.inter[1][0] ,
         \genblk1.inter[0][15] , \genblk1.inter[0][14] ,
         \genblk1.inter[0][13] , \genblk1.inter[0][12] ,
         \genblk1.inter[0][11] , \genblk1.inter[0][10] , \genblk1.inter[0][9] ,
         \genblk1.inter[0][8] , \genblk1.inter[0][7] , \genblk1.inter[0][6] ,
         \genblk1.inter[0][5] , \genblk1.inter[0][4] , \genblk1.inter[0][3] ,
         \genblk1.inter[0][2] , \genblk1.inter[0][1] , \genblk1.inter[0][0] ;

  recursive_add_layer_INPUT_SCALE2_WIDTH16_3 \genblk1.next_layer  ( .in({
        \genblk1.inter[1][15] , \genblk1.inter[1][14] , \genblk1.inter[1][13] , 
        \genblk1.inter[1][12] , \genblk1.inter[1][11] , \genblk1.inter[1][10] , 
        \genblk1.inter[1][9] , \genblk1.inter[1][8] , \genblk1.inter[1][7] , 
        \genblk1.inter[1][6] , \genblk1.inter[1][5] , \genblk1.inter[1][4] , 
        \genblk1.inter[1][3] , \genblk1.inter[1][2] , \genblk1.inter[1][1] , 
        \genblk1.inter[1][0] , \genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }), .out(out) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_3_DW01_add_4 add_64_G2 ( .A({
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] }), .B({\in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] }), .CI(1'b0), .SUM({\genblk1.inter[1][15] , \genblk1.inter[1][14] , 
        \genblk1.inter[1][13] , \genblk1.inter[1][12] , \genblk1.inter[1][11] , 
        \genblk1.inter[1][10] , \genblk1.inter[1][9] , \genblk1.inter[1][8] , 
        \genblk1.inter[1][7] , \genblk1.inter[1][6] , \genblk1.inter[1][5] , 
        \genblk1.inter[1][4] , \genblk1.inter[1][3] , \genblk1.inter[1][2] , 
        \genblk1.inter[1][1] , \genblk1.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_3_DW01_add_5 add_64 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM({\genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }) );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_3 ( .a({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , 
        \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , 
        \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , 
        \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , \x[1][7] , 
        \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , 
        \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , 
        \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \multout[3][15] , \multout[3][14] , \multout[3][13] ,
         \multout[3][12] , \multout[3][11] , \multout[3][10] , \multout[3][9] ,
         \multout[3][8] , \multout[3][7] , \multout[3][6] , \multout[3][5] ,
         \multout[3][4] , \multout[3][3] , \multout[3][2] , \multout[3][1] ,
         \multout[3][0] , \multout[2][15] , \multout[2][14] , \multout[2][13] ,
         \multout[2][12] , \multout[2][11] , \multout[2][10] , \multout[2][9] ,
         \multout[2][8] , \multout[2][7] , \multout[2][6] , \multout[2][5] ,
         \multout[2][4] , \multout[2][3] , \multout[2][2] , \multout[2][1] ,
         \multout[2][0] , \multout[1][15] , \multout[1][14] , \multout[1][13] ,
         \multout[1][12] , \multout[1][11] , \multout[1][10] , \multout[1][9] ,
         \multout[1][8] , \multout[1][7] , \multout[1][6] , \multout[1][5] ,
         \multout[1][4] , \multout[1][3] , \multout[1][2] , \multout[1][1] ,
         \multout[1][0] , \multout[0][15] , \multout[0][14] , \multout[0][13] ,
         \multout[0][12] , \multout[0][11] , \multout[0][10] , \multout[0][9] ,
         \multout[0][8] , \multout[0][7] , \multout[0][6] , \multout[0][5] ,
         \multout[0][4] , \multout[0][3] , \multout[0][2] , \multout[0][1] ,
         \multout[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_12 \genblk1[0].mult  ( .ia({\a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({\multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_11 \genblk1[1].mult  ( .ia({\a[1][7] , 
        \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , 
        \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , 
        \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({\multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_10 \genblk1[2].mult  ( .ia({\a[2][7] , 
        \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , \a[2][1] , 
        \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] , 
        \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({\multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_9 \genblk1[3].mult  ( .ia({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_3 add ( .in({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] , \multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] , \multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] , \multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n80, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100,
         n102, n103, n104, n108, n109, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n157, n158, n160, n161, n163, n164,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n245, n247, n248, n249, n250,
         n251, n252, n253, n255, n256, n258, n259, n260, n261, n262, n263,
         n264, n265, n273, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n332, n333,
         n334, n335, n336, n337;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n195), .B(n188), .CI(n182), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n189), .B(n177), .CI(n196), .CO(n144), .S(n145) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n199), .B(n192), .CO(n152), .S(n153) );
  NAND2_X1 U268 ( .A1(n249), .A2(n273), .ZN(n303) );
  NAND2_X1 U269 ( .A1(n249), .A2(n273), .ZN(n253) );
  CLKBUF_X3 U270 ( .A(n265), .Z(n314) );
  CLKBUF_X1 U271 ( .A(n263), .Z(n304) );
  OAI21_X1 U272 ( .B1(n61), .B2(n65), .A(n62), .ZN(n305) );
  OAI21_X1 U273 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  BUF_X1 U274 ( .A(n1), .Z(n335) );
  OR2_X1 U275 ( .A1(n137), .A2(n142), .ZN(n306) );
  NOR2_X2 U276 ( .A1(n64), .A2(n61), .ZN(n3) );
  OR2_X2 U277 ( .A1(n323), .A2(n324), .ZN(n307) );
  CLKBUF_X3 U278 ( .A(n245), .Z(n337) );
  OR2_X1 U279 ( .A1(n143), .A2(n146), .ZN(n308) );
  CLKBUF_X1 U280 ( .A(n263), .Z(n309) );
  BUF_X2 U281 ( .A(n327), .Z(n310) );
  XNOR2_X1 U282 ( .A(n263), .B(a[6]), .ZN(n327) );
  XNOR2_X1 U283 ( .A(n133), .B(n311), .ZN(n131) );
  XNOR2_X1 U284 ( .A(n138), .B(n135), .ZN(n311) );
  BUF_X1 U285 ( .A(n255), .Z(n332) );
  INV_X1 U286 ( .A(n64), .ZN(n103) );
  OR2_X1 U287 ( .A1(n201), .A2(n169), .ZN(n312) );
  BUF_X2 U288 ( .A(n264), .Z(n313) );
  XNOR2_X1 U289 ( .A(n261), .B(n164), .ZN(n249) );
  XOR2_X1 U290 ( .A(n190), .B(n197), .Z(n315) );
  XOR2_X1 U291 ( .A(n149), .B(n315), .Z(n147) );
  NAND2_X1 U292 ( .A1(n149), .A2(n190), .ZN(n316) );
  NAND2_X1 U293 ( .A1(n149), .A2(n197), .ZN(n317) );
  NAND2_X1 U294 ( .A1(n190), .A2(n197), .ZN(n318) );
  NAND3_X1 U295 ( .A1(n316), .A2(n317), .A3(n318), .ZN(n146) );
  CLKBUF_X1 U296 ( .A(n256), .Z(n336) );
  XNOR2_X1 U297 ( .A(n265), .B(a[2]), .ZN(n319) );
  NAND2_X1 U298 ( .A1(n133), .A2(n138), .ZN(n320) );
  NAND2_X1 U299 ( .A1(n133), .A2(n135), .ZN(n321) );
  NAND2_X1 U300 ( .A1(n138), .A2(n135), .ZN(n322) );
  NAND3_X1 U301 ( .A1(n320), .A2(n321), .A3(n322), .ZN(n130) );
  OR2_X2 U302 ( .A1(n323), .A2(n324), .ZN(n250) );
  XNOR2_X1 U303 ( .A(a[6]), .B(n262), .ZN(n323) );
  XOR2_X1 U304 ( .A(n263), .B(a[6]), .Z(n324) );
  NOR2_X1 U305 ( .A1(n131), .A2(n136), .ZN(n325) );
  NOR2_X1 U306 ( .A1(n131), .A2(n136), .ZN(n69) );
  XNOR2_X1 U307 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U308 ( .A1(n332), .A2(n247), .ZN(n326) );
  NOR2_X1 U309 ( .A1(n125), .A2(n130), .ZN(n64) );
  NAND2_X1 U310 ( .A1(n125), .A2(n130), .ZN(n65) );
  NOR2_X1 U311 ( .A1(n121), .A2(n124), .ZN(n61) );
  NOR2_X1 U312 ( .A1(n137), .A2(n142), .ZN(n72) );
  INV_X2 U313 ( .A(n164), .ZN(n273) );
  INV_X1 U314 ( .A(n30), .ZN(n28) );
  XNOR2_X1 U315 ( .A(n334), .B(n328), .ZN(product[9]) );
  AND2_X1 U316 ( .A1(n103), .A2(n65), .ZN(n328) );
  INV_X1 U317 ( .A(n31), .ZN(n29) );
  INV_X1 U318 ( .A(n18), .ZN(product[15]) );
  AOI21_X1 U319 ( .B1(n305), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U320 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  NAND2_X1 U321 ( .A1(n52), .A2(n32), .ZN(n30) );
  INV_X1 U322 ( .A(n305), .ZN(n58) );
  NAND2_X1 U323 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U324 ( .A(n61), .ZN(n102) );
  XNOR2_X1 U325 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U326 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U327 ( .A(n34), .ZN(n99) );
  XNOR2_X1 U328 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U329 ( .A1(n329), .A2(n94), .ZN(n16) );
  NAND2_X1 U330 ( .A1(n308), .A2(n77), .ZN(n12) );
  INV_X1 U331 ( .A(n82), .ZN(n80) );
  XNOR2_X1 U332 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U333 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U334 ( .A(n23), .ZN(n98) );
  NAND2_X1 U335 ( .A1(n306), .A2(n73), .ZN(n11) );
  XNOR2_X1 U336 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U337 ( .A1(n52), .A2(n51), .ZN(n7) );
  INV_X1 U338 ( .A(n50), .ZN(n52) );
  AOI21_X1 U339 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U340 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U341 ( .A1(n41), .A2(n34), .ZN(n32) );
  NAND2_X1 U342 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U343 ( .A(n41), .ZN(n100) );
  AOI21_X1 U344 ( .B1(n329), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U345 ( .A(n94), .ZN(n92) );
  XNOR2_X1 U346 ( .A(n13), .B(n83), .ZN(product[5]) );
  NAND2_X1 U347 ( .A1(n330), .A2(n82), .ZN(n13) );
  XNOR2_X1 U348 ( .A(n71), .B(n10), .ZN(product[8]) );
  NAND2_X1 U349 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U350 ( .A(n325), .ZN(n104) );
  OAI21_X1 U351 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  NOR2_X1 U352 ( .A1(n30), .A2(n23), .ZN(n21) );
  INV_X1 U353 ( .A(n51), .ZN(n53) );
  NOR2_X1 U354 ( .A1(n50), .A2(n41), .ZN(n39) );
  AOI21_X1 U355 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U356 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  NAND2_X1 U357 ( .A1(n131), .A2(n136), .ZN(n70) );
  XOR2_X1 U358 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U359 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U360 ( .A(n84), .ZN(n108) );
  NOR2_X1 U361 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U362 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U363 ( .A1(n187), .A2(n175), .ZN(n134) );
  XOR2_X1 U364 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U365 ( .A(n88), .ZN(n109) );
  NOR2_X1 U366 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U367 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U368 ( .A(n112), .ZN(n113) );
  NOR2_X1 U369 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U370 ( .A1(n170), .A2(n112), .ZN(n24) );
  OAI21_X1 U371 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  NAND2_X1 U372 ( .A1(n116), .A2(n115), .ZN(n44) );
  INV_X1 U373 ( .A(n97), .ZN(n95) );
  OR2_X1 U374 ( .A1(n200), .A2(n193), .ZN(n329) );
  NAND2_X1 U375 ( .A1(n117), .A2(n120), .ZN(n51) );
  NOR2_X1 U376 ( .A1(n143), .A2(n146), .ZN(n76) );
  INV_X1 U377 ( .A(n87), .ZN(n86) );
  NAND2_X1 U378 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U379 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U380 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U381 ( .A1(n147), .A2(n150), .ZN(n82) );
  NAND2_X1 U382 ( .A1(n143), .A2(n146), .ZN(n77) );
  OR2_X1 U383 ( .A1(n147), .A2(n150), .ZN(n330) );
  AND2_X1 U384 ( .A1(n337), .A2(n161), .ZN(n193) );
  AND2_X1 U385 ( .A1(n337), .A2(n158), .ZN(n185) );
  INV_X1 U386 ( .A(n157), .ZN(n178) );
  INV_X1 U387 ( .A(n118), .ZN(n119) );
  OR2_X1 U388 ( .A1(n337), .A2(n259), .ZN(n219) );
  NOR2_X1 U389 ( .A1(n151), .A2(n152), .ZN(n84) );
  BUF_X2 U390 ( .A(n255), .Z(n333) );
  AND2_X1 U391 ( .A1(n312), .A2(n97), .ZN(product[1]) );
  INV_X1 U392 ( .A(n163), .ZN(n194) );
  INV_X1 U393 ( .A(n128), .ZN(n129) );
  AND2_X1 U394 ( .A1(n337), .A2(n155), .ZN(n177) );
  NAND2_X1 U395 ( .A1(n151), .A2(n152), .ZN(n85) );
  INV_X1 U396 ( .A(n154), .ZN(n170) );
  OR2_X1 U397 ( .A1(n337), .A2(n258), .ZN(n210) );
  OR2_X1 U398 ( .A1(n337), .A2(n260), .ZN(n228) );
  OR2_X1 U399 ( .A1(n337), .A2(n261), .ZN(n237) );
  XNOR2_X1 U400 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U401 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U402 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U403 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U404 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U405 ( .A(b[4]), .B(n262), .ZN(n205) );
  NAND2_X1 U406 ( .A1(n247), .A2(n332), .ZN(n251) );
  XNOR2_X1 U407 ( .A(b[1]), .B(n262), .ZN(n208) );
  AND2_X1 U408 ( .A1(n337), .A2(n164), .ZN(product[0]) );
  XNOR2_X1 U409 ( .A(n262), .B(n337), .ZN(n209) );
  INV_X1 U410 ( .A(n262), .ZN(n258) );
  XNOR2_X1 U411 ( .A(n264), .B(a[4]), .ZN(n255) );
  OAI22_X1 U412 ( .A1(n303), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  OAI22_X1 U413 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  OAI22_X1 U414 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U415 ( .A1(n303), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U416 ( .A1(n229), .A2(n303), .B1(n229), .B2(n273), .ZN(n163) );
  OAI22_X1 U417 ( .A1(n303), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U418 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  INV_X1 U419 ( .A(n160), .ZN(n186) );
  NOR2_X1 U420 ( .A1(n153), .A2(n168), .ZN(n88) );
  BUF_X1 U421 ( .A(n1), .Z(n334) );
  NAND2_X1 U422 ( .A1(n200), .A2(n193), .ZN(n94) );
  OAI22_X1 U423 ( .A1(n303), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  XNOR2_X1 U424 ( .A(n265), .B(a[2]), .ZN(n256) );
  AOI21_X1 U425 ( .B1(n75), .B2(n67), .A(n68), .ZN(n1) );
  NAND2_X1 U426 ( .A1(n3), .A2(n21), .ZN(n19) );
  XNOR2_X1 U427 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U428 ( .A1(n3), .A2(n39), .ZN(n37) );
  INV_X1 U429 ( .A(n3), .ZN(n57) );
  NAND2_X1 U430 ( .A1(n3), .A2(n52), .ZN(n46) );
  OAI21_X1 U431 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NAND2_X1 U432 ( .A1(n109), .A2(n89), .ZN(n15) );
  AOI21_X1 U433 ( .B1(n330), .B2(n83), .A(n80), .ZN(n78) );
  OAI21_X1 U434 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  XOR2_X1 U435 ( .A(n12), .B(n78), .Z(product[6]) );
  OAI21_X1 U436 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  NOR2_X1 U437 ( .A1(n325), .A2(n72), .ZN(n67) );
  OAI21_X1 U438 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  XOR2_X1 U439 ( .A(n74), .B(n11), .Z(product[7]) );
  NAND2_X1 U440 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U441 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  NAND2_X1 U442 ( .A1(n3), .A2(n28), .ZN(n26) );
  AOI21_X1 U443 ( .B1(n305), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U444 ( .A(n75), .ZN(n74) );
  XNOR2_X1 U445 ( .A(b[2]), .B(n263), .ZN(n216) );
  XNOR2_X1 U446 ( .A(b[3]), .B(n263), .ZN(n215) );
  XNOR2_X1 U447 ( .A(b[4]), .B(n309), .ZN(n214) );
  XNOR2_X1 U448 ( .A(b[5]), .B(n304), .ZN(n213) );
  XNOR2_X1 U449 ( .A(b[7]), .B(n309), .ZN(n211) );
  XNOR2_X1 U450 ( .A(b[6]), .B(n263), .ZN(n212) );
  XNOR2_X1 U451 ( .A(n304), .B(n337), .ZN(n218) );
  INV_X1 U452 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U453 ( .A(b[1]), .B(n263), .ZN(n217) );
  XOR2_X1 U454 ( .A(n263), .B(a[4]), .Z(n247) );
  NAND2_X1 U455 ( .A1(n153), .A2(n168), .ZN(n89) );
  OAI22_X1 U456 ( .A1(n326), .A2(n217), .B1(n216), .B2(n333), .ZN(n183) );
  OAI22_X1 U457 ( .A1(n251), .A2(n216), .B1(n215), .B2(n333), .ZN(n182) );
  OAI22_X1 U458 ( .A1(n251), .A2(n212), .B1(n211), .B2(n333), .ZN(n118) );
  OAI22_X1 U459 ( .A1(n326), .A2(n215), .B1(n214), .B2(n333), .ZN(n181) );
  OAI22_X1 U460 ( .A1(n251), .A2(n214), .B1(n213), .B2(n333), .ZN(n180) );
  OAI22_X1 U461 ( .A1(n211), .A2(n326), .B1(n211), .B2(n333), .ZN(n157) );
  OAI22_X1 U462 ( .A1(n326), .A2(n213), .B1(n212), .B2(n333), .ZN(n179) );
  XNOR2_X1 U463 ( .A(b[5]), .B(n313), .ZN(n222) );
  INV_X1 U464 ( .A(n333), .ZN(n158) );
  OAI22_X1 U465 ( .A1(n251), .A2(n259), .B1(n219), .B2(n333), .ZN(n167) );
  OAI22_X1 U466 ( .A1(n251), .A2(n218), .B1(n217), .B2(n333), .ZN(n184) );
  XNOR2_X1 U467 ( .A(b[3]), .B(n313), .ZN(n224) );
  XNOR2_X1 U468 ( .A(b[4]), .B(n313), .ZN(n223) );
  XNOR2_X1 U469 ( .A(b[6]), .B(n313), .ZN(n221) );
  XNOR2_X1 U470 ( .A(b[2]), .B(n313), .ZN(n225) );
  INV_X1 U471 ( .A(n313), .ZN(n260) );
  XNOR2_X1 U472 ( .A(b[7]), .B(n313), .ZN(n220) );
  XNOR2_X1 U473 ( .A(n313), .B(n337), .ZN(n227) );
  XNOR2_X1 U474 ( .A(b[1]), .B(n313), .ZN(n226) );
  XOR2_X1 U475 ( .A(n264), .B(a[2]), .Z(n248) );
  OAI22_X1 U476 ( .A1(n202), .A2(n250), .B1(n202), .B2(n310), .ZN(n154) );
  OAI22_X1 U477 ( .A1(n307), .A2(n206), .B1(n205), .B2(n310), .ZN(n173) );
  OAI22_X1 U478 ( .A1(n307), .A2(n203), .B1(n202), .B2(n310), .ZN(n112) );
  OAI22_X1 U479 ( .A1(n250), .A2(n205), .B1(n204), .B2(n310), .ZN(n172) );
  OAI22_X1 U480 ( .A1(n250), .A2(n204), .B1(n203), .B2(n310), .ZN(n171) );
  OAI22_X1 U481 ( .A1(n307), .A2(n208), .B1(n207), .B2(n310), .ZN(n175) );
  OAI22_X1 U482 ( .A1(n250), .A2(n207), .B1(n206), .B2(n310), .ZN(n174) );
  INV_X1 U483 ( .A(n327), .ZN(n155) );
  OAI22_X1 U484 ( .A1(n307), .A2(n258), .B1(n210), .B2(n310), .ZN(n166) );
  OAI22_X1 U485 ( .A1(n250), .A2(n209), .B1(n208), .B2(n310), .ZN(n176) );
  OAI21_X1 U486 ( .B1(n334), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U487 ( .B1(n335), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U488 ( .B1(n335), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U489 ( .B1(n335), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U490 ( .B1(n334), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U491 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  OAI22_X1 U492 ( .A1(n252), .A2(n221), .B1(n220), .B2(n319), .ZN(n128) );
  OAI22_X1 U493 ( .A1(n220), .A2(n252), .B1(n220), .B2(n336), .ZN(n160) );
  OAI22_X1 U494 ( .A1(n252), .A2(n222), .B1(n221), .B2(n336), .ZN(n187) );
  OAI22_X1 U495 ( .A1(n252), .A2(n223), .B1(n222), .B2(n319), .ZN(n188) );
  OAI22_X1 U496 ( .A1(n252), .A2(n225), .B1(n224), .B2(n319), .ZN(n190) );
  OAI22_X1 U497 ( .A1(n252), .A2(n224), .B1(n223), .B2(n319), .ZN(n189) );
  OAI22_X1 U498 ( .A1(n252), .A2(n226), .B1(n225), .B2(n336), .ZN(n191) );
  OAI22_X1 U499 ( .A1(n252), .A2(n260), .B1(n228), .B2(n336), .ZN(n168) );
  XNOR2_X1 U500 ( .A(b[5]), .B(n314), .ZN(n231) );
  XNOR2_X1 U501 ( .A(b[6]), .B(n314), .ZN(n230) );
  XNOR2_X1 U502 ( .A(b[4]), .B(n314), .ZN(n232) );
  INV_X1 U503 ( .A(n319), .ZN(n161) );
  OAI22_X1 U504 ( .A1(n252), .A2(n227), .B1(n226), .B2(n336), .ZN(n192) );
  XNOR2_X1 U505 ( .A(b[7]), .B(n314), .ZN(n229) );
  NAND2_X2 U506 ( .A1(n248), .A2(n256), .ZN(n252) );
  XNOR2_X1 U507 ( .A(n314), .B(n337), .ZN(n236) );
  XNOR2_X1 U508 ( .A(b[3]), .B(n314), .ZN(n233) );
  XNOR2_X1 U509 ( .A(b[2]), .B(n314), .ZN(n234) );
  INV_X1 U510 ( .A(n265), .ZN(n261) );
  XNOR2_X1 U511 ( .A(b[1]), .B(n314), .ZN(n235) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50,
         n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102, n103,
         n104, n105, n108, n109, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n157, n158, n160, n161, n163, n164, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n245, n246, n247, n248, n249, n251,
         n252, n253, n254, n255, n256, n258, n259, n260, n261, n262, n263,
         n264, n265, n273, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n346, n347, n348, n349;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  CLKBUF_X1 U268 ( .A(n264), .Z(n303) );
  XOR2_X1 U269 ( .A(n194), .B(n181), .Z(n304) );
  XOR2_X1 U270 ( .A(n304), .B(n140), .Z(n133) );
  XOR2_X1 U271 ( .A(n138), .B(n135), .Z(n305) );
  XOR2_X1 U272 ( .A(n305), .B(n133), .Z(n131) );
  NAND2_X1 U273 ( .A1(n194), .A2(n181), .ZN(n306) );
  NAND2_X1 U274 ( .A1(n194), .A2(n140), .ZN(n307) );
  NAND2_X1 U275 ( .A1(n181), .A2(n140), .ZN(n308) );
  NAND3_X1 U276 ( .A1(n306), .A2(n307), .A3(n308), .ZN(n132) );
  NAND2_X1 U277 ( .A1(n138), .A2(n135), .ZN(n309) );
  NAND2_X1 U278 ( .A1(n138), .A2(n133), .ZN(n310) );
  NAND2_X1 U279 ( .A1(n135), .A2(n133), .ZN(n311) );
  NAND3_X1 U280 ( .A1(n309), .A2(n310), .A3(n311), .ZN(n130) );
  NAND2_X1 U281 ( .A1(n263), .A2(n313), .ZN(n314) );
  NAND2_X1 U282 ( .A1(n312), .A2(a[4]), .ZN(n315) );
  NAND2_X1 U283 ( .A1(n314), .A2(n315), .ZN(n247) );
  INV_X1 U284 ( .A(n263), .ZN(n312) );
  INV_X1 U285 ( .A(a[4]), .ZN(n313) );
  NOR2_X1 U286 ( .A1(n318), .A2(n72), .ZN(n316) );
  BUF_X2 U287 ( .A(n265), .Z(n320) );
  XNOR2_X1 U288 ( .A(n264), .B(a[4]), .ZN(n317) );
  NOR2_X1 U289 ( .A1(n131), .A2(n136), .ZN(n318) );
  NOR2_X1 U290 ( .A1(n131), .A2(n136), .ZN(n69) );
  CLKBUF_X1 U291 ( .A(n262), .Z(n319) );
  CLKBUF_X3 U292 ( .A(n256), .Z(n347) );
  OR2_X2 U293 ( .A1(n147), .A2(n150), .ZN(n343) );
  CLKBUF_X1 U294 ( .A(n263), .Z(n321) );
  XOR2_X1 U295 ( .A(a[6]), .B(n262), .Z(n322) );
  NOR2_X2 U296 ( .A1(n121), .A2(n124), .ZN(n61) );
  NOR2_X2 U297 ( .A1(n64), .A2(n61), .ZN(n3) );
  OR2_X1 U298 ( .A1(n143), .A2(n146), .ZN(n323) );
  BUF_X1 U299 ( .A(n256), .Z(n346) );
  OR2_X1 U300 ( .A1(n201), .A2(n169), .ZN(n324) );
  XNOR2_X1 U301 ( .A(n341), .B(n325), .ZN(product[9]) );
  AND2_X1 U302 ( .A1(n103), .A2(n65), .ZN(n325) );
  NAND2_X2 U303 ( .A1(n249), .A2(n273), .ZN(n253) );
  AOI21_X1 U304 ( .B1(n343), .B2(n83), .A(n334), .ZN(n326) );
  CLKBUF_X1 U305 ( .A(n340), .Z(n327) );
  NAND2_X1 U306 ( .A1(n248), .A2(n346), .ZN(n328) );
  NAND2_X1 U307 ( .A1(n248), .A2(n346), .ZN(n252) );
  NAND2_X1 U308 ( .A1(n246), .A2(n254), .ZN(n329) );
  NAND2_X1 U309 ( .A1(n322), .A2(n254), .ZN(n330) );
  OAI21_X2 U310 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  BUF_X2 U311 ( .A(n342), .Z(n331) );
  BUF_X1 U312 ( .A(n342), .Z(n332) );
  INV_X1 U313 ( .A(n334), .ZN(n82) );
  CLKBUF_X1 U314 ( .A(n83), .Z(n333) );
  AND2_X1 U315 ( .A1(n147), .A2(n150), .ZN(n334) );
  INV_X1 U316 ( .A(n260), .ZN(n335) );
  AOI21_X1 U317 ( .B1(n343), .B2(n83), .A(n334), .ZN(n78) );
  OAI21_X1 U318 ( .B1(n76), .B2(n326), .A(n77), .ZN(n336) );
  NAND2_X1 U319 ( .A1(n247), .A2(n317), .ZN(n337) );
  NAND2_X1 U320 ( .A1(n247), .A2(n317), .ZN(n338) );
  XOR2_X1 U321 ( .A(n339), .B(n326), .Z(product[6]) );
  NAND2_X1 U322 ( .A1(n323), .A2(n77), .ZN(n339) );
  BUF_X2 U323 ( .A(n245), .Z(n349) );
  INV_X2 U324 ( .A(n164), .ZN(n273) );
  AOI21_X1 U325 ( .B1(n336), .B2(n67), .A(n68), .ZN(n340) );
  AOI21_X1 U326 ( .B1(n316), .B2(n336), .A(n68), .ZN(n341) );
  XNOR2_X1 U327 ( .A(n263), .B(a[6]), .ZN(n342) );
  INV_X1 U328 ( .A(n30), .ZN(n28) );
  INV_X1 U329 ( .A(n64), .ZN(n103) );
  INV_X1 U330 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U331 ( .A1(n3), .A2(n21), .ZN(n19) );
  INV_X1 U332 ( .A(n31), .ZN(n29) );
  NAND2_X1 U333 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U334 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U335 ( .A1(n3), .A2(n39), .ZN(n37) );
  NAND2_X1 U336 ( .A1(n3), .A2(n28), .ZN(n26) );
  INV_X1 U337 ( .A(n3), .ZN(n57) );
  XNOR2_X1 U338 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U339 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U340 ( .A(n34), .ZN(n99) );
  XNOR2_X1 U341 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U342 ( .A1(n344), .A2(n94), .ZN(n16) );
  XNOR2_X1 U343 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U344 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U345 ( .A(n23), .ZN(n98) );
  XNOR2_X1 U346 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U347 ( .A1(n52), .A2(n51), .ZN(n7) );
  NAND2_X1 U348 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U349 ( .A(n318), .ZN(n104) );
  NAND2_X1 U350 ( .A1(n343), .A2(n82), .ZN(n13) );
  XNOR2_X1 U351 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U352 ( .A1(n102), .A2(n62), .ZN(n8) );
  XNOR2_X1 U353 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U354 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U355 ( .A(n41), .ZN(n100) );
  INV_X1 U356 ( .A(n50), .ZN(n52) );
  AOI21_X1 U357 ( .B1(n316), .B2(n336), .A(n68), .ZN(n1) );
  AOI21_X1 U358 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U359 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  OAI21_X1 U360 ( .B1(n76), .B2(n78), .A(n77), .ZN(n75) );
  NOR2_X1 U361 ( .A1(n125), .A2(n130), .ZN(n64) );
  XOR2_X1 U362 ( .A(n74), .B(n11), .Z(product[7]) );
  NAND2_X1 U363 ( .A1(n105), .A2(n73), .ZN(n11) );
  INV_X1 U364 ( .A(n72), .ZN(n105) );
  NOR2_X1 U365 ( .A1(n41), .A2(n34), .ZN(n32) );
  OAI21_X1 U366 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  AOI21_X1 U367 ( .B1(n344), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U368 ( .A(n94), .ZN(n92) );
  NOR2_X1 U369 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U370 ( .A1(n50), .A2(n41), .ZN(n39) );
  NAND2_X1 U371 ( .A1(n125), .A2(n130), .ZN(n65) );
  OAI21_X1 U372 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U373 ( .A(n51), .ZN(n53) );
  NAND2_X1 U374 ( .A1(n131), .A2(n136), .ZN(n70) );
  XOR2_X1 U375 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U376 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U377 ( .A(n84), .ZN(n108) );
  NOR2_X1 U378 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U379 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U380 ( .A1(n187), .A2(n175), .ZN(n134) );
  XOR2_X1 U381 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U382 ( .A(n88), .ZN(n109) );
  NOR2_X1 U383 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U384 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U385 ( .A(n112), .ZN(n113) );
  OAI21_X1 U386 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  NOR2_X1 U387 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U388 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U389 ( .A1(n116), .A2(n115), .ZN(n44) );
  INV_X1 U390 ( .A(n97), .ZN(n95) );
  NOR2_X1 U391 ( .A1(n137), .A2(n142), .ZN(n72) );
  OR2_X1 U392 ( .A1(n200), .A2(n193), .ZN(n344) );
  NOR2_X1 U393 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U394 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U395 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U396 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U397 ( .A1(n143), .A2(n146), .ZN(n77) );
  INV_X1 U398 ( .A(n87), .ZN(n86) );
  NAND2_X1 U399 ( .A1(n121), .A2(n124), .ZN(n62) );
  AND2_X1 U400 ( .A1(n349), .A2(n161), .ZN(n193) );
  AND2_X1 U401 ( .A1(n349), .A2(n158), .ZN(n185) );
  INV_X1 U402 ( .A(n157), .ZN(n178) );
  INV_X1 U403 ( .A(n118), .ZN(n119) );
  OR2_X1 U404 ( .A1(n349), .A2(n259), .ZN(n219) );
  NOR2_X1 U405 ( .A1(n153), .A2(n168), .ZN(n88) );
  AND2_X1 U406 ( .A1(n324), .A2(n97), .ZN(product[1]) );
  NOR2_X1 U407 ( .A1(n151), .A2(n152), .ZN(n84) );
  INV_X1 U408 ( .A(n163), .ZN(n194) );
  INV_X1 U409 ( .A(n128), .ZN(n129) );
  AND2_X1 U410 ( .A1(n349), .A2(n155), .ZN(n177) );
  INV_X1 U411 ( .A(n154), .ZN(n170) );
  NAND2_X1 U412 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U413 ( .A1(n349), .A2(n258), .ZN(n210) );
  XNOR2_X1 U414 ( .A(n263), .B(a[6]), .ZN(n254) );
  OR2_X1 U415 ( .A1(n349), .A2(n260), .ZN(n228) );
  OR2_X1 U416 ( .A1(n349), .A2(n261), .ZN(n237) );
  XNOR2_X1 U417 ( .A(b[7]), .B(n319), .ZN(n202) );
  XNOR2_X1 U418 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U419 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U420 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U421 ( .A(b[6]), .B(n262), .ZN(n203) );
  XOR2_X1 U422 ( .A(a[6]), .B(n262), .Z(n246) );
  NAND2_X1 U423 ( .A1(n247), .A2(n317), .ZN(n251) );
  XNOR2_X1 U424 ( .A(n262), .B(n349), .ZN(n209) );
  INV_X1 U425 ( .A(n262), .ZN(n258) );
  AND2_X1 U426 ( .A1(n349), .A2(n164), .ZN(product[0]) );
  NAND2_X1 U427 ( .A1(n109), .A2(n89), .ZN(n15) );
  OAI21_X1 U428 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  INV_X1 U429 ( .A(n160), .ZN(n186) );
  XNOR2_X1 U430 ( .A(n265), .B(a[2]), .ZN(n256) );
  BUF_X2 U431 ( .A(n255), .Z(n348) );
  XNOR2_X1 U432 ( .A(n13), .B(n333), .ZN(product[5]) );
  XNOR2_X1 U433 ( .A(n71), .B(n10), .ZN(product[8]) );
  XNOR2_X1 U434 ( .A(b[5]), .B(n335), .ZN(n222) );
  INV_X1 U435 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U436 ( .A(b[6]), .B(n303), .ZN(n221) );
  XNOR2_X1 U437 ( .A(b[3]), .B(n264), .ZN(n224) );
  XNOR2_X1 U438 ( .A(b[7]), .B(n264), .ZN(n220) );
  XNOR2_X1 U439 ( .A(b[4]), .B(n264), .ZN(n223) );
  XNOR2_X1 U440 ( .A(n303), .B(n349), .ZN(n227) );
  XOR2_X1 U441 ( .A(n264), .B(a[2]), .Z(n248) );
  XNOR2_X1 U442 ( .A(n264), .B(a[4]), .ZN(n255) );
  AOI21_X1 U443 ( .B1(n2), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U444 ( .B1(n2), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U445 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  INV_X1 U446 ( .A(n2), .ZN(n58) );
  INV_X1 U447 ( .A(n61), .ZN(n102) );
  AOI21_X1 U448 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  OAI21_X1 U449 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  NOR2_X1 U450 ( .A1(n318), .A2(n72), .ZN(n67) );
  OAI21_X1 U451 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  NAND2_X1 U452 ( .A1(n200), .A2(n193), .ZN(n94) );
  XNOR2_X1 U453 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U454 ( .A(b[2]), .B(n303), .ZN(n225) );
  INV_X1 U455 ( .A(n75), .ZN(n74) );
  XNOR2_X1 U456 ( .A(b[1]), .B(n262), .ZN(n208) );
  XNOR2_X1 U457 ( .A(b[1]), .B(n264), .ZN(n226) );
  OAI22_X1 U458 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  OAI22_X1 U459 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  NAND2_X1 U460 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U461 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U462 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U463 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  OAI22_X1 U464 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U465 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OAI22_X1 U466 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OAI22_X1 U467 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OAI22_X1 U468 ( .A1(n338), .A2(n217), .B1(n216), .B2(n348), .ZN(n183) );
  OAI22_X1 U469 ( .A1(n337), .A2(n212), .B1(n211), .B2(n348), .ZN(n118) );
  OAI22_X1 U470 ( .A1(n337), .A2(n216), .B1(n215), .B2(n348), .ZN(n182) );
  OAI22_X1 U471 ( .A1(n338), .A2(n215), .B1(n214), .B2(n348), .ZN(n181) );
  OAI22_X1 U472 ( .A1(n211), .A2(n338), .B1(n211), .B2(n348), .ZN(n157) );
  OAI22_X1 U473 ( .A1(n338), .A2(n214), .B1(n213), .B2(n348), .ZN(n180) );
  OAI22_X1 U474 ( .A1(n337), .A2(n213), .B1(n212), .B2(n348), .ZN(n179) );
  OAI22_X1 U475 ( .A1(n251), .A2(n259), .B1(n219), .B2(n348), .ZN(n167) );
  OAI22_X1 U476 ( .A1(n251), .A2(n218), .B1(n217), .B2(n348), .ZN(n184) );
  INV_X1 U477 ( .A(n348), .ZN(n158) );
  NAND2_X1 U478 ( .A1(n153), .A2(n168), .ZN(n89) );
  XNOR2_X1 U479 ( .A(b[5]), .B(n320), .ZN(n231) );
  XNOR2_X1 U480 ( .A(b[6]), .B(n320), .ZN(n230) );
  XNOR2_X1 U481 ( .A(b[4]), .B(n320), .ZN(n232) );
  XNOR2_X1 U482 ( .A(b[7]), .B(n265), .ZN(n229) );
  XNOR2_X1 U483 ( .A(n320), .B(n349), .ZN(n236) );
  XNOR2_X1 U484 ( .A(b[2]), .B(n320), .ZN(n234) );
  XNOR2_X1 U485 ( .A(b[3]), .B(n320), .ZN(n233) );
  XNOR2_X1 U486 ( .A(b[1]), .B(n320), .ZN(n235) );
  INV_X1 U487 ( .A(n265), .ZN(n261) );
  XOR2_X1 U488 ( .A(n265), .B(n164), .Z(n249) );
  OAI22_X1 U489 ( .A1(n202), .A2(n329), .B1(n202), .B2(n331), .ZN(n154) );
  OAI22_X1 U490 ( .A1(n329), .A2(n206), .B1(n205), .B2(n331), .ZN(n173) );
  OAI22_X1 U491 ( .A1(n330), .A2(n203), .B1(n202), .B2(n332), .ZN(n112) );
  OAI22_X1 U492 ( .A1(n329), .A2(n205), .B1(n204), .B2(n331), .ZN(n172) );
  OAI22_X1 U493 ( .A1(n330), .A2(n204), .B1(n203), .B2(n332), .ZN(n171) );
  OAI22_X1 U494 ( .A1(n330), .A2(n208), .B1(n207), .B2(n332), .ZN(n175) );
  OAI22_X1 U495 ( .A1(n329), .A2(n207), .B1(n206), .B2(n331), .ZN(n174) );
  INV_X1 U496 ( .A(n342), .ZN(n155) );
  OAI22_X1 U497 ( .A1(n329), .A2(n258), .B1(n210), .B2(n332), .ZN(n166) );
  OAI22_X1 U498 ( .A1(n330), .A2(n209), .B1(n208), .B2(n331), .ZN(n176) );
  XNOR2_X1 U499 ( .A(b[2]), .B(n321), .ZN(n216) );
  XNOR2_X1 U500 ( .A(b[3]), .B(n263), .ZN(n215) );
  XNOR2_X1 U501 ( .A(b[4]), .B(n263), .ZN(n214) );
  XNOR2_X1 U502 ( .A(b[7]), .B(n321), .ZN(n211) );
  XNOR2_X1 U503 ( .A(b[5]), .B(n321), .ZN(n213) );
  XNOR2_X1 U504 ( .A(b[6]), .B(n263), .ZN(n212) );
  XNOR2_X1 U505 ( .A(n263), .B(n349), .ZN(n218) );
  INV_X1 U506 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U507 ( .A(b[1]), .B(n263), .ZN(n217) );
  OAI21_X1 U508 ( .B1(n327), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U509 ( .B1(n341), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U510 ( .B1(n340), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U511 ( .B1(n341), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U512 ( .B1(n340), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U513 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  OAI22_X1 U514 ( .A1(n252), .A2(n221), .B1(n220), .B2(n347), .ZN(n128) );
  OAI22_X1 U515 ( .A1(n220), .A2(n328), .B1(n220), .B2(n347), .ZN(n160) );
  OAI22_X1 U516 ( .A1(n252), .A2(n222), .B1(n221), .B2(n347), .ZN(n187) );
  OAI22_X1 U517 ( .A1(n252), .A2(n224), .B1(n223), .B2(n347), .ZN(n189) );
  OAI22_X1 U518 ( .A1(n328), .A2(n225), .B1(n224), .B2(n347), .ZN(n190) );
  OAI22_X1 U519 ( .A1(n328), .A2(n223), .B1(n222), .B2(n347), .ZN(n188) );
  OAI22_X1 U520 ( .A1(n328), .A2(n260), .B1(n228), .B2(n347), .ZN(n168) );
  OAI22_X1 U521 ( .A1(n328), .A2(n226), .B1(n225), .B2(n347), .ZN(n191) );
  OAI22_X1 U522 ( .A1(n252), .A2(n227), .B1(n226), .B2(n347), .ZN(n192) );
  INV_X1 U523 ( .A(n347), .ZN(n161) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50, n51, n52,
         n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n92, n94, n95, n97, n98, n99, n100, n102, n103, n105, n108,
         n109, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n157, n158, n160, n161, n163, n164, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n258, n259, n260, n261, n262, n263, n264, n265,
         n273, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n345, n346,
         n347, n348, n349, n350, n351, n352;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n320), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n129), .B(n180), .CI(n174), .CO(n126), .S(n127) );
  FA_X1 U136 ( .A(n138), .B(n135), .CI(n133), .CO(n130), .S(n131) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n167), .B(n184), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n199), .B(n192), .CO(n152), .S(n153) );
  INV_X1 U268 ( .A(n262), .ZN(n303) );
  INV_X2 U269 ( .A(n303), .ZN(n304) );
  NOR2_X1 U270 ( .A1(n121), .A2(n124), .ZN(n305) );
  NOR2_X1 U271 ( .A1(n121), .A2(n124), .ZN(n306) );
  NOR2_X1 U272 ( .A1(n121), .A2(n124), .ZN(n61) );
  INV_X1 U273 ( .A(n103), .ZN(n307) );
  AOI21_X1 U274 ( .B1(n342), .B2(n83), .A(n331), .ZN(n308) );
  AOI21_X1 U275 ( .B1(n342), .B2(n83), .A(n331), .ZN(n78) );
  CLKBUF_X1 U276 ( .A(n70), .Z(n309) );
  OAI21_X1 U277 ( .B1(n76), .B2(n308), .A(n77), .ZN(n310) );
  CLKBUF_X1 U278 ( .A(n304), .Z(n311) );
  CLKBUF_X1 U279 ( .A(n332), .Z(n312) );
  BUF_X2 U280 ( .A(n265), .Z(n351) );
  CLKBUF_X1 U281 ( .A(n83), .Z(n313) );
  BUF_X2 U282 ( .A(n255), .Z(n347) );
  BUF_X2 U283 ( .A(n255), .Z(n346) );
  OR2_X1 U284 ( .A1(n147), .A2(n150), .ZN(n342) );
  NOR2_X1 U285 ( .A1(n137), .A2(n142), .ZN(n72) );
  NOR2_X1 U286 ( .A1(n125), .A2(n130), .ZN(n64) );
  CLKBUF_X1 U287 ( .A(n264), .Z(n314) );
  BUF_X1 U288 ( .A(n256), .Z(n348) );
  CLKBUF_X1 U289 ( .A(n264), .Z(n315) );
  BUF_X1 U290 ( .A(n1), .Z(n316) );
  OR2_X1 U291 ( .A1(n143), .A2(n146), .ZN(n317) );
  XNOR2_X1 U292 ( .A(n264), .B(a[4]), .ZN(n318) );
  BUF_X2 U293 ( .A(n263), .Z(n333) );
  BUF_X1 U294 ( .A(n254), .Z(n345) );
  INV_X1 U295 ( .A(n261), .ZN(n319) );
  OAI22_X1 U296 ( .A1(n332), .A2(n221), .B1(n220), .B2(n349), .ZN(n320) );
  CLKBUF_X1 U297 ( .A(n256), .Z(n349) );
  CLKBUF_X1 U298 ( .A(n256), .Z(n350) );
  OAI22_X1 U299 ( .A1(n332), .A2(n221), .B1(n220), .B2(n349), .ZN(n128) );
  BUF_X2 U300 ( .A(n245), .Z(n352) );
  INV_X1 U301 ( .A(n72), .ZN(n105) );
  OR2_X1 U302 ( .A1(n323), .A2(n136), .ZN(n321) );
  OR2_X1 U303 ( .A1(n201), .A2(n169), .ZN(n322) );
  FA_X1 U304 ( .A(n138), .B(n135), .CI(n133), .S(n323) );
  OAI21_X1 U305 ( .B1(n305), .B2(n65), .A(n62), .ZN(n324) );
  OAI21_X1 U306 ( .B1(n306), .B2(n65), .A(n62), .ZN(n325) );
  OAI21_X1 U307 ( .B1(n306), .B2(n65), .A(n62), .ZN(n2) );
  AOI21_X1 U308 ( .B1(n67), .B2(n310), .A(n68), .ZN(n336) );
  NOR2_X2 U309 ( .A1(n64), .A2(n61), .ZN(n3) );
  XNOR2_X1 U310 ( .A(n263), .B(a[6]), .ZN(n326) );
  CLKBUF_X1 U311 ( .A(n263), .Z(n327) );
  INV_X1 U312 ( .A(n331), .ZN(n82) );
  AND2_X1 U313 ( .A1(n147), .A2(n150), .ZN(n331) );
  NOR2_X1 U314 ( .A1(n131), .A2(n136), .ZN(n328) );
  NOR2_X1 U315 ( .A1(n131), .A2(n136), .ZN(n69) );
  XNOR2_X1 U316 ( .A(n336), .B(n329), .ZN(product[9]) );
  AND2_X1 U317 ( .A1(n103), .A2(n65), .ZN(n329) );
  CLKBUF_X1 U318 ( .A(n251), .Z(n330) );
  NAND2_X1 U319 ( .A1(n318), .A2(n247), .ZN(n251) );
  NAND2_X1 U320 ( .A1(n248), .A2(n348), .ZN(n332) );
  NAND2_X1 U321 ( .A1(n248), .A2(n348), .ZN(n252) );
  CLKBUF_X1 U322 ( .A(n336), .Z(n334) );
  CLKBUF_X1 U323 ( .A(n308), .Z(n335) );
  AOI21_X1 U324 ( .B1(n67), .B2(n310), .A(n68), .ZN(n1) );
  INV_X1 U325 ( .A(n250), .ZN(n337) );
  INV_X1 U326 ( .A(n337), .ZN(n338) );
  XNOR2_X1 U327 ( .A(n339), .B(n313), .ZN(product[5]) );
  NAND2_X1 U328 ( .A1(n342), .A2(n82), .ZN(n339) );
  XOR2_X1 U329 ( .A(n74), .B(n340), .Z(product[7]) );
  NAND2_X1 U330 ( .A1(n105), .A2(n73), .ZN(n340) );
  XOR2_X1 U331 ( .A(n341), .B(n335), .Z(product[6]) );
  NAND2_X1 U332 ( .A1(n317), .A2(n77), .ZN(n341) );
  NOR2_X1 U333 ( .A1(n143), .A2(n146), .ZN(n76) );
  INV_X1 U334 ( .A(n30), .ZN(n28) );
  INV_X1 U335 ( .A(n64), .ZN(n103) );
  AOI21_X1 U336 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  AOI21_X1 U337 ( .B1(n325), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U338 ( .A(n31), .ZN(n29) );
  NAND2_X1 U339 ( .A1(n52), .A2(n32), .ZN(n30) );
  INV_X1 U340 ( .A(n75), .ZN(n74) );
  INV_X1 U341 ( .A(n324), .ZN(n58) );
  INV_X1 U342 ( .A(n18), .ZN(product[15]) );
  AOI21_X1 U343 ( .B1(n324), .B2(n21), .A(n22), .ZN(n20) );
  NAND2_X1 U344 ( .A1(n3), .A2(n21), .ZN(n19) );
  NAND2_X1 U345 ( .A1(n3), .A2(n39), .ZN(n37) );
  NAND2_X1 U346 ( .A1(n3), .A2(n28), .ZN(n26) );
  NAND2_X1 U347 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U348 ( .A(n305), .ZN(n102) );
  XNOR2_X1 U349 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U350 ( .A1(n343), .A2(n94), .ZN(n16) );
  NAND2_X1 U351 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U352 ( .A(n41), .ZN(n100) );
  NAND2_X1 U353 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U354 ( .A(n23), .ZN(n98) );
  XNOR2_X1 U355 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U356 ( .A1(n52), .A2(n51), .ZN(n7) );
  INV_X1 U357 ( .A(n3), .ZN(n57) );
  XNOR2_X1 U358 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U359 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U360 ( .A(n34), .ZN(n99) );
  NAND2_X1 U361 ( .A1(n321), .A2(n309), .ZN(n10) );
  OAI21_X1 U362 ( .B1(n76), .B2(n78), .A(n77), .ZN(n75) );
  INV_X1 U363 ( .A(n50), .ZN(n52) );
  AOI21_X1 U364 ( .B1(n343), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U365 ( .A(n94), .ZN(n92) );
  AOI21_X1 U366 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U367 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U368 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U369 ( .A1(n50), .A2(n41), .ZN(n39) );
  NOR2_X1 U370 ( .A1(n41), .A2(n34), .ZN(n32) );
  OAI21_X1 U371 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U372 ( .A(n51), .ZN(n53) );
  NAND2_X1 U373 ( .A1(n125), .A2(n130), .ZN(n65) );
  AOI21_X1 U374 ( .B1(n325), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U375 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  NAND2_X1 U376 ( .A1(n323), .A2(n136), .ZN(n70) );
  XOR2_X1 U377 ( .A(n15), .B(n90), .Z(product[3]) );
  NAND2_X1 U378 ( .A1(n109), .A2(n89), .ZN(n15) );
  INV_X1 U379 ( .A(n88), .ZN(n109) );
  NOR2_X1 U380 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U381 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U382 ( .A1(n187), .A2(n175), .ZN(n134) );
  XOR2_X1 U383 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U384 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U385 ( .A(n84), .ZN(n108) );
  OR2_X1 U386 ( .A1(n200), .A2(n193), .ZN(n343) );
  NOR2_X1 U387 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U388 ( .A1(n114), .A2(n113), .ZN(n34) );
  OAI21_X1 U389 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  INV_X1 U390 ( .A(n112), .ZN(n113) );
  NOR2_X1 U391 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U392 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U393 ( .A1(n116), .A2(n115), .ZN(n44) );
  INV_X1 U394 ( .A(n97), .ZN(n95) );
  NAND2_X1 U395 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U396 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U397 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U398 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U399 ( .A1(n143), .A2(n146), .ZN(n77) );
  INV_X1 U400 ( .A(n87), .ZN(n86) );
  OAI21_X1 U401 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  AND2_X1 U402 ( .A1(n352), .A2(n161), .ZN(n193) );
  INV_X1 U403 ( .A(n157), .ZN(n178) );
  INV_X1 U404 ( .A(n118), .ZN(n119) );
  AND2_X1 U405 ( .A1(n352), .A2(n158), .ZN(n185) );
  OAI22_X1 U406 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U407 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OR2_X1 U408 ( .A1(n352), .A2(n259), .ZN(n219) );
  OAI22_X1 U409 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  NOR2_X1 U410 ( .A1(n153), .A2(n168), .ZN(n88) );
  AND2_X1 U411 ( .A1(n322), .A2(n97), .ZN(product[1]) );
  NOR2_X1 U412 ( .A1(n151), .A2(n152), .ZN(n84) );
  INV_X1 U413 ( .A(n160), .ZN(n186) );
  INV_X1 U414 ( .A(n128), .ZN(n129) );
  AND2_X1 U415 ( .A1(n352), .A2(n155), .ZN(n177) );
  OAI22_X1 U416 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U417 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  INV_X1 U418 ( .A(n154), .ZN(n170) );
  NAND2_X1 U419 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U420 ( .A1(n352), .A2(n258), .ZN(n210) );
  INV_X1 U421 ( .A(n163), .ZN(n194) );
  OAI22_X1 U422 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  OR2_X1 U423 ( .A1(n352), .A2(n260), .ZN(n228) );
  OR2_X1 U424 ( .A1(n352), .A2(n261), .ZN(n237) );
  NAND2_X1 U425 ( .A1(n246), .A2(n254), .ZN(n250) );
  AND2_X1 U426 ( .A1(n245), .A2(n164), .ZN(product[0]) );
  OAI22_X1 U427 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  XNOR2_X1 U428 ( .A(n263), .B(a[6]), .ZN(n254) );
  XNOR2_X1 U429 ( .A(n264), .B(a[4]), .ZN(n255) );
  NAND2_X1 U430 ( .A1(n200), .A2(n193), .ZN(n94) );
  XNOR2_X1 U431 ( .A(n265), .B(a[2]), .ZN(n256) );
  XNOR2_X1 U432 ( .A(n63), .B(n8), .ZN(product[10]) );
  OAI21_X1 U433 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  NOR2_X1 U434 ( .A1(n328), .A2(n72), .ZN(n67) );
  NAND2_X1 U435 ( .A1(n3), .A2(n52), .ZN(n46) );
  XNOR2_X1 U436 ( .A(n45), .B(n6), .ZN(product[12]) );
  XNOR2_X1 U437 ( .A(n304), .B(b[4]), .ZN(n205) );
  XNOR2_X1 U438 ( .A(b[7]), .B(n311), .ZN(n202) );
  XNOR2_X1 U439 ( .A(b[5]), .B(n304), .ZN(n204) );
  XNOR2_X1 U440 ( .A(b[6]), .B(n304), .ZN(n203) );
  XNOR2_X1 U441 ( .A(b[2]), .B(n304), .ZN(n207) );
  XNOR2_X1 U442 ( .A(n262), .B(b[3]), .ZN(n206) );
  XNOR2_X1 U443 ( .A(n262), .B(n352), .ZN(n209) );
  INV_X1 U444 ( .A(n262), .ZN(n258) );
  XNOR2_X1 U445 ( .A(b[1]), .B(n262), .ZN(n208) );
  XOR2_X1 U446 ( .A(n262), .B(a[6]), .Z(n246) );
  NAND2_X1 U447 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U448 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OAI22_X1 U449 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  NAND2_X2 U450 ( .A1(n249), .A2(n273), .ZN(n253) );
  XNOR2_X1 U451 ( .A(n25), .B(n4), .ZN(product[14]) );
  OAI22_X1 U452 ( .A1(n202), .A2(n338), .B1(n202), .B2(n345), .ZN(n154) );
  OAI22_X1 U453 ( .A1(n338), .A2(n206), .B1(n205), .B2(n326), .ZN(n173) );
  OAI22_X1 U454 ( .A1(n338), .A2(n203), .B1(n202), .B2(n326), .ZN(n112) );
  OAI22_X1 U455 ( .A1(n338), .A2(n205), .B1(n204), .B2(n345), .ZN(n172) );
  OAI22_X1 U456 ( .A1(n338), .A2(n208), .B1(n207), .B2(n326), .ZN(n175) );
  OAI22_X1 U457 ( .A1(n338), .A2(n204), .B1(n203), .B2(n345), .ZN(n171) );
  OAI22_X1 U458 ( .A1(n338), .A2(n207), .B1(n206), .B2(n345), .ZN(n174) );
  OAI22_X1 U459 ( .A1(n250), .A2(n258), .B1(n210), .B2(n326), .ZN(n166) );
  OAI22_X1 U460 ( .A1(n250), .A2(n209), .B1(n208), .B2(n345), .ZN(n176) );
  XNOR2_X1 U461 ( .A(b[2]), .B(n327), .ZN(n216) );
  XNOR2_X1 U462 ( .A(b[3]), .B(n333), .ZN(n215) );
  XNOR2_X1 U463 ( .A(b[4]), .B(n327), .ZN(n214) );
  INV_X1 U464 ( .A(n326), .ZN(n155) );
  XNOR2_X1 U465 ( .A(n333), .B(n352), .ZN(n218) );
  XNOR2_X1 U466 ( .A(b[6]), .B(n333), .ZN(n212) );
  XNOR2_X1 U467 ( .A(b[5]), .B(n333), .ZN(n213) );
  XNOR2_X1 U468 ( .A(b[7]), .B(n333), .ZN(n211) );
  XNOR2_X1 U469 ( .A(b[1]), .B(n327), .ZN(n217) );
  INV_X1 U470 ( .A(n333), .ZN(n259) );
  XOR2_X1 U471 ( .A(n263), .B(a[4]), .Z(n247) );
  XNOR2_X1 U472 ( .A(n71), .B(n10), .ZN(product[8]) );
  OAI21_X1 U473 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  OAI22_X1 U474 ( .A1(n330), .A2(n217), .B1(n216), .B2(n346), .ZN(n183) );
  OAI22_X1 U475 ( .A1(n251), .A2(n215), .B1(n214), .B2(n347), .ZN(n181) );
  OAI22_X1 U476 ( .A1(n330), .A2(n212), .B1(n211), .B2(n347), .ZN(n118) );
  OAI22_X1 U477 ( .A1(n251), .A2(n216), .B1(n215), .B2(n346), .ZN(n182) );
  OAI22_X1 U478 ( .A1(n211), .A2(n330), .B1(n211), .B2(n346), .ZN(n157) );
  OAI22_X1 U479 ( .A1(n251), .A2(n214), .B1(n213), .B2(n346), .ZN(n180) );
  OAI22_X1 U480 ( .A1(n251), .A2(n213), .B1(n212), .B2(n347), .ZN(n179) );
  OAI22_X1 U481 ( .A1(n251), .A2(n259), .B1(n219), .B2(n347), .ZN(n167) );
  OAI22_X1 U482 ( .A1(n251), .A2(n218), .B1(n217), .B2(n346), .ZN(n184) );
  INV_X1 U483 ( .A(n347), .ZN(n158) );
  NAND2_X1 U484 ( .A1(n153), .A2(n168), .ZN(n89) );
  XNOR2_X1 U485 ( .A(b[5]), .B(n315), .ZN(n222) );
  XNOR2_X1 U486 ( .A(b[3]), .B(n314), .ZN(n224) );
  XNOR2_X1 U487 ( .A(b[4]), .B(n264), .ZN(n223) );
  INV_X1 U488 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U489 ( .A(b[6]), .B(n314), .ZN(n221) );
  XNOR2_X1 U490 ( .A(b[2]), .B(n315), .ZN(n225) );
  XNOR2_X1 U491 ( .A(b[7]), .B(n264), .ZN(n220) );
  XNOR2_X1 U492 ( .A(n264), .B(n352), .ZN(n227) );
  XNOR2_X1 U493 ( .A(b[1]), .B(n264), .ZN(n226) );
  XOR2_X1 U494 ( .A(n264), .B(a[2]), .Z(n248) );
  OAI21_X1 U495 ( .B1(n334), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U496 ( .B1(n316), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U497 ( .B1(n316), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U498 ( .B1(n336), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U499 ( .B1(n336), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U500 ( .B1(n1), .B2(n307), .A(n65), .ZN(n63) );
  OAI22_X1 U501 ( .A1(n220), .A2(n332), .B1(n220), .B2(n350), .ZN(n160) );
  OAI22_X1 U502 ( .A1(n252), .A2(n222), .B1(n221), .B2(n350), .ZN(n187) );
  OAI22_X1 U503 ( .A1(n252), .A2(n224), .B1(n223), .B2(n350), .ZN(n189) );
  OAI22_X1 U504 ( .A1(n312), .A2(n225), .B1(n224), .B2(n349), .ZN(n190) );
  OAI22_X1 U505 ( .A1(n332), .A2(n223), .B1(n222), .B2(n350), .ZN(n188) );
  OAI22_X1 U506 ( .A1(n312), .A2(n260), .B1(n228), .B2(n349), .ZN(n168) );
  OAI22_X1 U507 ( .A1(n332), .A2(n226), .B1(n225), .B2(n349), .ZN(n191) );
  XNOR2_X1 U508 ( .A(b[5]), .B(n351), .ZN(n231) );
  XNOR2_X1 U509 ( .A(b[6]), .B(n351), .ZN(n230) );
  INV_X1 U510 ( .A(n349), .ZN(n161) );
  XNOR2_X1 U511 ( .A(b[4]), .B(n351), .ZN(n232) );
  OAI22_X1 U512 ( .A1(n252), .A2(n227), .B1(n226), .B2(n350), .ZN(n192) );
  XNOR2_X1 U513 ( .A(b[7]), .B(n319), .ZN(n229) );
  XNOR2_X1 U514 ( .A(n351), .B(n352), .ZN(n236) );
  XNOR2_X1 U515 ( .A(b[3]), .B(n351), .ZN(n233) );
  XNOR2_X1 U516 ( .A(b[2]), .B(n319), .ZN(n234) );
  INV_X1 U517 ( .A(n265), .ZN(n261) );
  XNOR2_X1 U518 ( .A(b[1]), .B(n351), .ZN(n235) );
  XOR2_X1 U519 ( .A(n265), .B(n164), .Z(n249) );
  INV_X2 U520 ( .A(n164), .ZN(n273) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102,
         n103, n104, n105, n108, n109, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n157, n160, n161, n163, n164, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n245, n246, n248, n250, n251, n252,
         n253, n254, n256, n258, n259, n260, n261, n262, n263, n264, n265,
         n273, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n341, n342, n343;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  NAND2_X1 U268 ( .A1(a[6]), .A2(n304), .ZN(n305) );
  NAND2_X1 U269 ( .A1(n303), .A2(n262), .ZN(n306) );
  NAND2_X1 U270 ( .A1(n305), .A2(n306), .ZN(n246) );
  INV_X1 U271 ( .A(a[6]), .ZN(n303) );
  INV_X1 U272 ( .A(n262), .ZN(n304) );
  OR2_X2 U273 ( .A1(n331), .A2(n330), .ZN(n307) );
  OR2_X2 U274 ( .A1(n308), .A2(n164), .ZN(n253) );
  XNOR2_X1 U275 ( .A(n265), .B(n164), .ZN(n308) );
  BUF_X1 U276 ( .A(n83), .Z(n309) );
  INV_X1 U277 ( .A(n164), .ZN(n273) );
  OAI21_X1 U278 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  CLKBUF_X1 U279 ( .A(n263), .Z(n310) );
  CLKBUF_X1 U280 ( .A(n263), .Z(n311) );
  BUF_X1 U281 ( .A(n263), .Z(n314) );
  CLKBUF_X1 U282 ( .A(n317), .Z(n312) );
  CLKBUF_X1 U283 ( .A(n264), .Z(n319) );
  BUF_X1 U284 ( .A(n264), .Z(n320) );
  XNOR2_X1 U285 ( .A(n336), .B(n313), .ZN(product[9]) );
  AND2_X1 U286 ( .A1(n103), .A2(n65), .ZN(n313) );
  BUF_X2 U287 ( .A(n254), .Z(n341) );
  BUF_X1 U288 ( .A(n263), .Z(n322) );
  BUF_X2 U289 ( .A(n265), .Z(n315) );
  AND2_X1 U290 ( .A1(n147), .A2(n150), .ZN(n317) );
  INV_X1 U291 ( .A(n317), .ZN(n82) );
  CLKBUF_X1 U292 ( .A(n338), .Z(n316) );
  BUF_X1 U293 ( .A(n1), .Z(n335) );
  OR2_X1 U294 ( .A1(n201), .A2(n169), .ZN(n318) );
  XNOR2_X1 U295 ( .A(n133), .B(n321), .ZN(n131) );
  XNOR2_X1 U296 ( .A(n135), .B(n138), .ZN(n321) );
  NOR2_X2 U297 ( .A1(n121), .A2(n124), .ZN(n61) );
  OR2_X1 U298 ( .A1(n143), .A2(n146), .ZN(n323) );
  NOR2_X2 U299 ( .A1(n64), .A2(n61), .ZN(n3) );
  AOI21_X1 U300 ( .B1(n309), .B2(n316), .A(n312), .ZN(n324) );
  XNOR2_X2 U301 ( .A(n264), .B(a[4]), .ZN(n337) );
  CLKBUF_X1 U302 ( .A(n265), .Z(n325) );
  OAI21_X2 U303 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  AND2_X1 U304 ( .A1(n246), .A2(n341), .ZN(n326) );
  NAND2_X1 U305 ( .A1(n133), .A2(n135), .ZN(n327) );
  NAND2_X1 U306 ( .A1(n133), .A2(n138), .ZN(n328) );
  NAND2_X1 U307 ( .A1(n135), .A2(n138), .ZN(n329) );
  NAND3_X1 U308 ( .A1(n327), .A2(n328), .A3(n329), .ZN(n130) );
  BUF_X1 U309 ( .A(n1), .Z(n336) );
  OR2_X2 U310 ( .A1(n331), .A2(n330), .ZN(n251) );
  XNOR2_X1 U311 ( .A(n314), .B(a[4]), .ZN(n330) );
  XOR2_X1 U312 ( .A(n264), .B(a[4]), .Z(n331) );
  XNOR2_X1 U313 ( .A(n265), .B(a[2]), .ZN(n332) );
  INV_X1 U314 ( .A(n326), .ZN(n333) );
  NAND2_X1 U315 ( .A1(n246), .A2(n254), .ZN(n250) );
  NOR2_X1 U316 ( .A1(n131), .A2(n136), .ZN(n334) );
  AOI21_X1 U317 ( .B1(n75), .B2(n67), .A(n68), .ZN(n1) );
  NOR2_X1 U318 ( .A1(n131), .A2(n136), .ZN(n69) );
  OR2_X1 U319 ( .A1(n147), .A2(n150), .ZN(n338) );
  CLKBUF_X3 U320 ( .A(n245), .Z(n343) );
  INV_X1 U321 ( .A(n30), .ZN(n28) );
  INV_X1 U322 ( .A(n64), .ZN(n103) );
  INV_X1 U323 ( .A(n18), .ZN(product[15]) );
  INV_X1 U324 ( .A(n31), .ZN(n29) );
  NAND2_X1 U325 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U326 ( .A1(n323), .A2(n77), .ZN(n12) );
  XNOR2_X1 U327 ( .A(n13), .B(n309), .ZN(product[5]) );
  NAND2_X1 U328 ( .A1(n316), .A2(n82), .ZN(n13) );
  NAND2_X1 U329 ( .A1(n105), .A2(n73), .ZN(n11) );
  INV_X1 U330 ( .A(n72), .ZN(n105) );
  XNOR2_X1 U331 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U332 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U333 ( .A(n61), .ZN(n102) );
  XNOR2_X1 U334 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U335 ( .A1(n52), .A2(n51), .ZN(n7) );
  XNOR2_X1 U336 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U337 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U338 ( .A(n34), .ZN(n99) );
  XNOR2_X1 U339 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U340 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U341 ( .A(n23), .ZN(n98) );
  AOI21_X1 U342 ( .B1(n339), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U343 ( .A(n94), .ZN(n92) );
  AOI21_X1 U344 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U345 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U346 ( .A1(n125), .A2(n130), .ZN(n64) );
  NOR2_X1 U347 ( .A1(n41), .A2(n34), .ZN(n32) );
  OAI21_X1 U348 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  NAND2_X1 U349 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U350 ( .A(n41), .ZN(n100) );
  INV_X1 U351 ( .A(n50), .ZN(n52) );
  XNOR2_X1 U352 ( .A(n71), .B(n10), .ZN(product[8]) );
  NAND2_X1 U353 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U354 ( .A(n334), .ZN(n104) );
  NAND2_X1 U355 ( .A1(n125), .A2(n130), .ZN(n65) );
  OAI21_X1 U356 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U357 ( .A(n51), .ZN(n53) );
  NOR2_X1 U358 ( .A1(n30), .A2(n23), .ZN(n21) );
  NAND2_X1 U359 ( .A1(n131), .A2(n136), .ZN(n70) );
  NOR2_X1 U360 ( .A1(n50), .A2(n41), .ZN(n39) );
  XNOR2_X1 U361 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U362 ( .A1(n339), .A2(n94), .ZN(n16) );
  NOR2_X1 U363 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U364 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U365 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U366 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U367 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U368 ( .A(n112), .ZN(n113) );
  NOR2_X1 U369 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U370 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U371 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U372 ( .A1(n137), .A2(n142), .ZN(n72) );
  INV_X1 U373 ( .A(n97), .ZN(n95) );
  XOR2_X1 U374 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U375 ( .A(n88), .ZN(n109) );
  OR2_X1 U376 ( .A1(n200), .A2(n193), .ZN(n339) );
  NAND2_X1 U377 ( .A1(n117), .A2(n120), .ZN(n51) );
  NOR2_X1 U378 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U379 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U380 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U381 ( .A1(n143), .A2(n146), .ZN(n77) );
  NAND2_X1 U382 ( .A1(n121), .A2(n124), .ZN(n62) );
  INV_X1 U383 ( .A(n87), .ZN(n86) );
  OAI21_X1 U384 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  AND2_X1 U385 ( .A1(n343), .A2(n161), .ZN(n193) );
  NAND2_X1 U386 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U387 ( .A(n84), .ZN(n108) );
  INV_X1 U388 ( .A(n157), .ZN(n178) );
  OAI22_X1 U389 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  AND2_X1 U390 ( .A1(n343), .A2(n331), .ZN(n185) );
  INV_X1 U391 ( .A(n118), .ZN(n119) );
  OAI22_X1 U392 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OR2_X1 U393 ( .A1(n343), .A2(n259), .ZN(n219) );
  NOR2_X1 U394 ( .A1(n153), .A2(n168), .ZN(n88) );
  AND2_X1 U395 ( .A1(n318), .A2(n97), .ZN(product[1]) );
  NOR2_X1 U396 ( .A1(n151), .A2(n152), .ZN(n84) );
  INV_X1 U397 ( .A(n163), .ZN(n194) );
  OAI22_X1 U398 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  INV_X1 U399 ( .A(n160), .ZN(n186) );
  INV_X1 U400 ( .A(n128), .ZN(n129) );
  OAI22_X1 U401 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  INV_X1 U402 ( .A(n154), .ZN(n170) );
  NAND2_X1 U403 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U404 ( .A1(n343), .A2(n258), .ZN(n210) );
  OAI22_X1 U405 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  AND2_X1 U406 ( .A1(n343), .A2(n155), .ZN(n177) );
  OR2_X1 U407 ( .A1(n343), .A2(n260), .ZN(n228) );
  OAI22_X1 U408 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OAI22_X1 U409 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OR2_X1 U410 ( .A1(n343), .A2(n261), .ZN(n237) );
  XNOR2_X1 U411 ( .A(n310), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U412 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U413 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U414 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U415 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U416 ( .A(n322), .B(b[7]), .ZN(n211) );
  XNOR2_X1 U417 ( .A(n262), .B(n343), .ZN(n209) );
  XNOR2_X1 U418 ( .A(n310), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U419 ( .A(n311), .B(b[6]), .ZN(n212) );
  INV_X1 U420 ( .A(n262), .ZN(n258) );
  AND2_X1 U421 ( .A1(n343), .A2(n164), .ZN(product[0]) );
  XNOR2_X1 U422 ( .A(n322), .B(n343), .ZN(n218) );
  INV_X1 U423 ( .A(n322), .ZN(n259) );
  XOR2_X1 U424 ( .A(n12), .B(n324), .Z(product[6]) );
  XNOR2_X1 U425 ( .A(n263), .B(a[6]), .ZN(n254) );
  BUF_X2 U426 ( .A(n256), .Z(n342) );
  XNOR2_X1 U427 ( .A(n265), .B(a[2]), .ZN(n256) );
  NAND2_X1 U428 ( .A1(n153), .A2(n168), .ZN(n89) );
  AOI21_X1 U429 ( .B1(n2), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U430 ( .B1(n2), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U431 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U432 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  INV_X1 U433 ( .A(n2), .ZN(n58) );
  XOR2_X1 U434 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U435 ( .A1(n3), .A2(n21), .ZN(n19) );
  NAND2_X1 U436 ( .A1(n3), .A2(n28), .ZN(n26) );
  INV_X1 U437 ( .A(n3), .ZN(n57) );
  NAND2_X1 U438 ( .A1(n3), .A2(n39), .ZN(n37) );
  NAND2_X1 U439 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U440 ( .A1(n200), .A2(n193), .ZN(n94) );
  XOR2_X1 U441 ( .A(n74), .B(n11), .Z(product[7]) );
  OAI21_X1 U442 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  INV_X1 U443 ( .A(n75), .ZN(n74) );
  OAI21_X1 U444 ( .B1(n76), .B2(n78), .A(n77), .ZN(n75) );
  AOI21_X1 U445 ( .B1(n83), .B2(n338), .A(n317), .ZN(n78) );
  OAI21_X1 U446 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  NOR2_X1 U447 ( .A1(n334), .A2(n72), .ZN(n67) );
  NAND2_X1 U448 ( .A1(n109), .A2(n89), .ZN(n15) );
  OAI22_X1 U449 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  XNOR2_X1 U450 ( .A(n310), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U451 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U452 ( .A(n311), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U453 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U454 ( .A(b[1]), .B(n262), .ZN(n208) );
  XNOR2_X1 U455 ( .A(n311), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U456 ( .A(n45), .B(n6), .ZN(product[12]) );
  OAI22_X1 U457 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  NAND2_X1 U458 ( .A1(n201), .A2(n169), .ZN(n97) );
  XNOR2_X1 U459 ( .A(n315), .B(b[5]), .ZN(n231) );
  XNOR2_X1 U460 ( .A(n315), .B(b[6]), .ZN(n230) );
  XNOR2_X1 U461 ( .A(n325), .B(b[4]), .ZN(n232) );
  XNOR2_X1 U462 ( .A(n315), .B(b[7]), .ZN(n229) );
  XNOR2_X1 U463 ( .A(n315), .B(b[2]), .ZN(n234) );
  XNOR2_X1 U464 ( .A(n315), .B(b[3]), .ZN(n233) );
  XNOR2_X1 U465 ( .A(n325), .B(n343), .ZN(n236) );
  XNOR2_X1 U466 ( .A(n315), .B(b[1]), .ZN(n235) );
  INV_X1 U467 ( .A(n265), .ZN(n261) );
  OAI21_X1 U468 ( .B1(n335), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U469 ( .B1(n335), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U470 ( .B1(n336), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U471 ( .B1(n336), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U472 ( .B1(n335), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U473 ( .B1(n64), .B2(n1), .A(n65), .ZN(n63) );
  OAI22_X1 U474 ( .A1(n202), .A2(n333), .B1(n202), .B2(n341), .ZN(n154) );
  OAI22_X1 U475 ( .A1(n333), .A2(n206), .B1(n341), .B2(n205), .ZN(n173) );
  OAI22_X1 U476 ( .A1(n333), .A2(n203), .B1(n341), .B2(n202), .ZN(n112) );
  OAI22_X1 U477 ( .A1(n333), .A2(n205), .B1(n341), .B2(n204), .ZN(n172) );
  OAI22_X1 U478 ( .A1(n333), .A2(n204), .B1(n341), .B2(n203), .ZN(n171) );
  OAI22_X1 U479 ( .A1(n250), .A2(n207), .B1(n341), .B2(n206), .ZN(n174) );
  OAI22_X1 U480 ( .A1(n250), .A2(n208), .B1(n341), .B2(n207), .ZN(n175) );
  INV_X1 U481 ( .A(n341), .ZN(n155) );
  OAI22_X1 U482 ( .A1(n250), .A2(n258), .B1(n210), .B2(n341), .ZN(n166) );
  OAI22_X1 U483 ( .A1(n250), .A2(n209), .B1(n341), .B2(n208), .ZN(n176) );
  OAI22_X1 U484 ( .A1(n251), .A2(n217), .B1(n216), .B2(n337), .ZN(n183) );
  OAI22_X1 U485 ( .A1(n307), .A2(n212), .B1(n211), .B2(n337), .ZN(n118) );
  OAI22_X1 U486 ( .A1(n211), .A2(n251), .B1(n211), .B2(n337), .ZN(n157) );
  OAI22_X1 U487 ( .A1(n307), .A2(n213), .B1(n212), .B2(n337), .ZN(n179) );
  OAI22_X1 U488 ( .A1(n251), .A2(n214), .B1(n213), .B2(n337), .ZN(n180) );
  OAI22_X1 U489 ( .A1(n251), .A2(n216), .B1(n215), .B2(n337), .ZN(n182) );
  OAI22_X1 U490 ( .A1(n307), .A2(n215), .B1(n214), .B2(n337), .ZN(n181) );
  XNOR2_X1 U491 ( .A(n319), .B(b[4]), .ZN(n223) );
  XNOR2_X1 U492 ( .A(n320), .B(b[6]), .ZN(n221) );
  XNOR2_X1 U493 ( .A(n320), .B(b[5]), .ZN(n222) );
  XNOR2_X1 U494 ( .A(n319), .B(b[3]), .ZN(n224) );
  OAI22_X1 U495 ( .A1(n307), .A2(n259), .B1(n219), .B2(n337), .ZN(n167) );
  OAI22_X1 U496 ( .A1(n251), .A2(n218), .B1(n217), .B2(n337), .ZN(n184) );
  INV_X1 U497 ( .A(n319), .ZN(n260) );
  XNOR2_X1 U498 ( .A(n320), .B(b[7]), .ZN(n220) );
  XNOR2_X1 U499 ( .A(n320), .B(b[2]), .ZN(n225) );
  XNOR2_X1 U500 ( .A(n319), .B(n343), .ZN(n227) );
  XNOR2_X1 U501 ( .A(n320), .B(b[1]), .ZN(n226) );
  XOR2_X1 U502 ( .A(n264), .B(a[2]), .Z(n248) );
  OAI22_X1 U503 ( .A1(n252), .A2(n222), .B1(n221), .B2(n342), .ZN(n187) );
  OAI22_X1 U504 ( .A1(n252), .A2(n224), .B1(n223), .B2(n332), .ZN(n189) );
  OAI22_X1 U505 ( .A1(n252), .A2(n221), .B1(n220), .B2(n332), .ZN(n128) );
  OAI22_X1 U506 ( .A1(n252), .A2(n225), .B1(n224), .B2(n342), .ZN(n190) );
  OAI22_X1 U507 ( .A1(n252), .A2(n223), .B1(n222), .B2(n332), .ZN(n188) );
  OAI22_X1 U508 ( .A1(n252), .A2(n260), .B1(n228), .B2(n332), .ZN(n168) );
  OAI22_X1 U509 ( .A1(n220), .A2(n252), .B1(n220), .B2(n342), .ZN(n160) );
  OAI22_X1 U510 ( .A1(n252), .A2(n226), .B1(n225), .B2(n342), .ZN(n191) );
  OAI22_X1 U511 ( .A1(n252), .A2(n227), .B1(n226), .B2(n332), .ZN(n192) );
  INV_X1 U512 ( .A(n342), .ZN(n161) );
  NAND2_X2 U513 ( .A1(n248), .A2(n256), .ZN(n252) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_2_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n20, n21, n22, n26, n27, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n51, n52, n54, n56,
         n57, n58, n60, n62, n63, n64, n65, n66, n68, n70, n71, n72, n73, n74,
         n76, n78, n79, n80, n81, n82, n84, n86, n87, n89, n93, n94, n95, n99,
         n101, n103, n160, n161, n162, n163, n164, n165, n166, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185;

  AND2_X1 U125 ( .A1(A[14]), .A2(B[14]), .ZN(n160) );
  INV_X4 U126 ( .A(n160), .ZN(n26) );
  CLKBUF_X1 U127 ( .A(n182), .Z(n161) );
  AOI21_X1 U128 ( .B1(n71), .B2(n181), .A(n68), .ZN(n162) );
  XNOR2_X1 U129 ( .A(n1), .B(n163), .ZN(SUM[12]) );
  AND2_X1 U130 ( .A1(n93), .A2(n174), .ZN(n163) );
  CLKBUF_X1 U131 ( .A(A[13]), .Z(n164) );
  CLKBUF_X1 U132 ( .A(n33), .Z(n166) );
  OR2_X1 U133 ( .A1(n172), .A2(n35), .ZN(n165) );
  CLKBUF_X1 U134 ( .A(B[13]), .Z(n171) );
  AOI21_X1 U135 ( .B1(n71), .B2(n181), .A(n68), .ZN(n66) );
  AND2_X1 U136 ( .A1(n169), .A2(n89), .ZN(SUM[0]) );
  OR2_X1 U137 ( .A1(B[7]), .A2(A[7]), .ZN(n168) );
  OR2_X1 U138 ( .A1(B[0]), .A2(A[0]), .ZN(n169) );
  XNOR2_X1 U139 ( .A(n44), .B(n170), .ZN(SUM[10]) );
  AND2_X1 U140 ( .A1(n95), .A2(n43), .ZN(n170) );
  OR2_X2 U141 ( .A1(B[14]), .A2(A[14]), .ZN(n182) );
  NOR2_X1 U142 ( .A1(B[13]), .A2(A[13]), .ZN(n172) );
  AOI21_X1 U143 ( .B1(n37), .B2(n45), .A(n38), .ZN(n173) );
  AOI21_X1 U144 ( .B1(n37), .B2(n45), .A(n38), .ZN(n1) );
  CLKBUF_X1 U145 ( .A(n36), .Z(n174) );
  NOR2_X1 U146 ( .A1(A[13]), .A2(B[13]), .ZN(n32) );
  OR2_X1 U147 ( .A1(A[9]), .A2(B[9]), .ZN(n175) );
  OR2_X1 U148 ( .A1(A[9]), .A2(B[9]), .ZN(n179) );
  OR2_X1 U149 ( .A1(n171), .A2(n164), .ZN(n176) );
  INV_X1 U150 ( .A(n177), .ZN(n51) );
  AND2_X1 U151 ( .A1(A[9]), .A2(B[9]), .ZN(n177) );
  NOR2_X1 U152 ( .A1(A[11]), .A2(B[11]), .ZN(n178) );
  NOR2_X1 U153 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  INV_X1 U154 ( .A(n58), .ZN(n57) );
  INV_X1 U155 ( .A(n62), .ZN(n60) );
  INV_X1 U156 ( .A(n42), .ZN(n95) );
  INV_X1 U157 ( .A(n35), .ZN(n93) );
  NAND2_X1 U158 ( .A1(n176), .A2(n166), .ZN(n4) );
  AOI21_X1 U159 ( .B1(n180), .B2(n57), .A(n54), .ZN(n52) );
  XOR2_X1 U160 ( .A(n11), .B(n162), .Z(SUM[6]) );
  NAND2_X1 U161 ( .A1(n99), .A2(n65), .ZN(n11) );
  INV_X1 U162 ( .A(n64), .ZN(n99) );
  XNOR2_X1 U163 ( .A(n9), .B(n57), .ZN(SUM[8]) );
  NAND2_X1 U164 ( .A1(n94), .A2(n40), .ZN(n6) );
  INV_X1 U165 ( .A(n178), .ZN(n94) );
  XNOR2_X1 U166 ( .A(n12), .B(n71), .ZN(SUM[5]) );
  NAND2_X1 U167 ( .A1(n181), .A2(n70), .ZN(n12) );
  INV_X1 U168 ( .A(n70), .ZN(n68) );
  NAND2_X1 U169 ( .A1(n168), .A2(n62), .ZN(n10) );
  OAI21_X1 U170 ( .B1(n72), .B2(n74), .A(n73), .ZN(n71) );
  AOI21_X1 U171 ( .B1(n184), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U172 ( .A(n78), .ZN(n76) );
  NAND2_X1 U173 ( .A1(B[10]), .A2(A[10]), .ZN(n43) );
  OR2_X1 U174 ( .A1(B[8]), .A2(A[8]), .ZN(n180) );
  NOR2_X1 U175 ( .A1(B[6]), .A2(A[6]), .ZN(n64) );
  OR2_X1 U176 ( .A1(B[5]), .A2(A[5]), .ZN(n181) );
  NAND2_X1 U177 ( .A1(B[6]), .A2(A[6]), .ZN(n65) );
  NAND2_X1 U178 ( .A1(n101), .A2(n73), .ZN(n13) );
  INV_X1 U179 ( .A(n72), .ZN(n101) );
  XNOR2_X1 U180 ( .A(n14), .B(n79), .ZN(SUM[3]) );
  NAND2_X1 U181 ( .A1(n184), .A2(n78), .ZN(n14) );
  OR2_X1 U182 ( .A1(B[15]), .A2(A[15]), .ZN(n183) );
  OAI21_X1 U183 ( .B1(n82), .B2(n80), .A(n81), .ZN(n79) );
  NAND2_X1 U184 ( .A1(B[4]), .A2(A[4]), .ZN(n73) );
  NOR2_X1 U185 ( .A1(B[4]), .A2(A[4]), .ZN(n72) );
  XOR2_X1 U186 ( .A(n15), .B(n82), .Z(SUM[2]) );
  NAND2_X1 U187 ( .A1(n103), .A2(n81), .ZN(n15) );
  INV_X1 U188 ( .A(n80), .ZN(n103) );
  OR2_X1 U189 ( .A1(B[3]), .A2(A[3]), .ZN(n184) );
  AOI21_X1 U190 ( .B1(n185), .B2(n87), .A(n84), .ZN(n82) );
  INV_X1 U191 ( .A(n86), .ZN(n84) );
  NOR2_X1 U192 ( .A1(B[2]), .A2(A[2]), .ZN(n80) );
  NAND2_X1 U193 ( .A1(B[2]), .A2(A[2]), .ZN(n81) );
  XNOR2_X1 U194 ( .A(n16), .B(n87), .ZN(SUM[1]) );
  NAND2_X1 U195 ( .A1(n185), .A2(n86), .ZN(n16) );
  OR2_X1 U196 ( .A1(B[1]), .A2(A[1]), .ZN(n185) );
  INV_X1 U197 ( .A(n89), .ZN(n87) );
  NAND2_X1 U198 ( .A1(B[1]), .A2(A[1]), .ZN(n86) );
  NAND2_X1 U199 ( .A1(B[0]), .A2(A[0]), .ZN(n89) );
  XNOR2_X1 U200 ( .A(n41), .B(n6), .ZN(SUM[11]) );
  XOR2_X1 U201 ( .A(n8), .B(n52), .Z(SUM[9]) );
  NAND2_X1 U202 ( .A1(n161), .A2(n26), .ZN(n3) );
  NAND2_X1 U203 ( .A1(n180), .A2(n56), .ZN(n9) );
  INV_X1 U204 ( .A(n56), .ZN(n54) );
  XNOR2_X1 U205 ( .A(n10), .B(n63), .ZN(SUM[7]) );
  NAND2_X1 U206 ( .A1(B[5]), .A2(A[5]), .ZN(n70) );
  OAI21_X1 U207 ( .B1(n64), .B2(n66), .A(n65), .ZN(n63) );
  NAND2_X1 U208 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  XOR2_X1 U209 ( .A(n13), .B(n74), .Z(SUM[4]) );
  NAND2_X1 U210 ( .A1(B[3]), .A2(A[3]), .ZN(n78) );
  NAND2_X1 U211 ( .A1(B[8]), .A2(A[8]), .ZN(n56) );
  NAND2_X1 U212 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  OAI21_X1 U213 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U214 ( .A1(A[13]), .A2(B[13]), .ZN(n33) );
  NAND2_X1 U215 ( .A1(n183), .A2(n19), .ZN(n2) );
  AOI21_X1 U216 ( .B1(n168), .B2(n63), .A(n60), .ZN(n58) );
  NOR2_X1 U217 ( .A1(A[12]), .A2(B[12]), .ZN(n35) );
  NAND2_X1 U218 ( .A1(B[12]), .A2(A[12]), .ZN(n36) );
  NOR2_X1 U219 ( .A1(B[10]), .A2(A[10]), .ZN(n42) );
  OAI21_X1 U220 ( .B1(n44), .B2(n42), .A(n43), .ZN(n41) );
  INV_X1 U221 ( .A(n45), .ZN(n44) );
  AOI21_X1 U222 ( .B1(n179), .B2(n54), .A(n177), .ZN(n47) );
  XNOR2_X1 U223 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U224 ( .A1(A[11]), .A2(B[11]), .ZN(n40) );
  XNOR2_X1 U225 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  OAI21_X1 U226 ( .B1(n46), .B2(n58), .A(n47), .ZN(n45) );
  INV_X1 U227 ( .A(n31), .ZN(n29) );
  AOI21_X1 U228 ( .B1(n31), .B2(n182), .A(n160), .ZN(n22) );
  NAND2_X1 U229 ( .A1(n30), .A2(n182), .ZN(n21) );
  OAI21_X1 U230 ( .B1(n39), .B2(n43), .A(n40), .ZN(n38) );
  NOR2_X1 U231 ( .A1(n178), .A2(n42), .ZN(n37) );
  NOR2_X1 U232 ( .A1(n172), .A2(n35), .ZN(n30) );
  XNOR2_X1 U233 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  OAI21_X1 U234 ( .B1(n173), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U235 ( .B1(n1), .B2(n165), .A(n29), .ZN(n27) );
  OAI21_X1 U236 ( .B1(n173), .B2(n35), .A(n174), .ZN(n34) );
  NAND2_X1 U237 ( .A1(n175), .A2(n51), .ZN(n8) );
  NAND2_X1 U238 ( .A1(n175), .A2(n180), .ZN(n46) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_2 ( .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;


  recursive_add_layer_INPUT_SCALE2_WIDTH16_2_DW01_add_2 add_56 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM(out) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_2_DW01_add_4 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n10, n12, n13, n14, n15, n16, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n36, n37, n38,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n59, n60, n62, n64, n65, n66, n68, n70, n71, n72, n73, n74,
         n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89, n91, n93, n94,
         n97, n98, n102, n104, n106, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189;

  CLKBUF_X1 U127 ( .A(B[11]), .Z(n162) );
  BUF_X1 U128 ( .A(n66), .Z(n163) );
  CLKBUF_X1 U129 ( .A(A[12]), .Z(n164) );
  CLKBUF_X1 U130 ( .A(n38), .Z(n165) );
  OR2_X1 U131 ( .A1(n42), .A2(n39), .ZN(n166) );
  CLKBUF_X1 U132 ( .A(n43), .Z(n167) );
  OR2_X1 U133 ( .A1(n162), .A2(A[11]), .ZN(n168) );
  NOR2_X1 U134 ( .A1(A[12]), .A2(B[12]), .ZN(n169) );
  OR2_X1 U135 ( .A1(n164), .A2(B[12]), .ZN(n170) );
  INV_X1 U136 ( .A(n166), .ZN(n171) );
  OR2_X1 U137 ( .A1(B[7]), .A2(A[7]), .ZN(n172) );
  AND2_X1 U138 ( .A1(n182), .A2(n91), .ZN(SUM[0]) );
  OAI21_X1 U139 ( .B1(n54), .B2(n163), .A(n175), .ZN(n174) );
  AOI21_X1 U140 ( .B1(n185), .B2(n62), .A(n178), .ZN(n175) );
  XNOR2_X1 U141 ( .A(n174), .B(n176), .ZN(SUM[9]) );
  NAND2_X1 U142 ( .A1(n98), .A2(n51), .ZN(n176) );
  NOR2_X1 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n177) );
  NOR2_X1 U144 ( .A1(A[10]), .A2(B[10]), .ZN(n47) );
  INV_X1 U145 ( .A(n178), .ZN(n59) );
  AND2_X1 U146 ( .A1(A[8]), .A2(B[8]), .ZN(n178) );
  OR2_X2 U147 ( .A1(A[8]), .A2(B[8]), .ZN(n185) );
  XNOR2_X1 U148 ( .A(n49), .B(n179), .ZN(SUM[10]) );
  NAND2_X1 U149 ( .A1(n97), .A2(n48), .ZN(n179) );
  NOR2_X1 U150 ( .A1(B[9]), .A2(A[9]), .ZN(n50) );
  AOI21_X1 U151 ( .B1(n53), .B2(n45), .A(n46), .ZN(n180) );
  AOI21_X1 U152 ( .B1(n53), .B2(n45), .A(n46), .ZN(n1) );
  AOI21_X1 U153 ( .B1(n186), .B2(n71), .A(n68), .ZN(n66) );
  XOR2_X1 U154 ( .A(n181), .B(n71), .Z(SUM[6]) );
  AND2_X1 U155 ( .A1(n186), .A2(n70), .ZN(n181) );
  OR2_X1 U156 ( .A1(B[6]), .A2(A[6]), .ZN(n186) );
  OR2_X1 U157 ( .A1(B[0]), .A2(A[0]), .ZN(n182) );
  INV_X1 U158 ( .A(n50), .ZN(n98) );
  INV_X1 U159 ( .A(n66), .ZN(n65) );
  NAND2_X1 U160 ( .A1(n37), .A2(n94), .ZN(n28) );
  NAND2_X1 U161 ( .A1(n171), .A2(n23), .ZN(n21) );
  NAND2_X1 U162 ( .A1(n94), .A2(n33), .ZN(n4) );
  OAI21_X1 U163 ( .B1(n54), .B2(n163), .A(n55), .ZN(n53) );
  NAND2_X1 U164 ( .A1(n172), .A2(n64), .ZN(n10) );
  NOR2_X1 U165 ( .A1(n42), .A2(n39), .ZN(n37) );
  XNOR2_X1 U166 ( .A(n60), .B(n183), .ZN(SUM[8]) );
  AND2_X1 U167 ( .A1(n185), .A2(n59), .ZN(n183) );
  OAI21_X1 U168 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  XOR2_X1 U169 ( .A(n12), .B(n74), .Z(SUM[5]) );
  NAND2_X1 U170 ( .A1(n102), .A2(n73), .ZN(n12) );
  INV_X1 U171 ( .A(n72), .ZN(n102) );
  INV_X1 U172 ( .A(n33), .ZN(n31) );
  NAND2_X1 U173 ( .A1(n170), .A2(n40), .ZN(n5) );
  NAND2_X1 U174 ( .A1(n93), .A2(n26), .ZN(n3) );
  INV_X1 U175 ( .A(n25), .ZN(n93) );
  NAND2_X1 U176 ( .A1(n184), .A2(n19), .ZN(n2) );
  NAND2_X1 U177 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  INV_X1 U178 ( .A(n70), .ZN(n68) );
  INV_X1 U179 ( .A(n32), .ZN(n94) );
  NOR2_X1 U180 ( .A1(n32), .A2(n25), .ZN(n23) );
  NAND2_X1 U181 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  OAI21_X1 U182 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  INV_X1 U183 ( .A(n64), .ZN(n62) );
  OR2_X1 U184 ( .A1(B[15]), .A2(A[15]), .ZN(n184) );
  NAND2_X1 U185 ( .A1(n188), .A2(n78), .ZN(n13) );
  NOR2_X1 U186 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  INV_X1 U187 ( .A(n78), .ZN(n76) );
  NOR2_X1 U188 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  NOR2_X1 U189 ( .A1(B[11]), .A2(A[11]), .ZN(n42) );
  NOR2_X1 U190 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  XOR2_X1 U191 ( .A(n14), .B(n82), .Z(SUM[3]) );
  INV_X1 U192 ( .A(n80), .ZN(n104) );
  NAND2_X1 U193 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  NOR2_X1 U194 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND2_X1 U195 ( .A1(A[13]), .A2(B[13]), .ZN(n33) );
  NAND2_X1 U196 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U197 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  NAND2_X1 U198 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
  OR2_X1 U199 ( .A1(B[2]), .A2(A[2]), .ZN(n187) );
  XNOR2_X1 U200 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U201 ( .A1(n187), .A2(n86), .ZN(n15) );
  AOI21_X1 U202 ( .B1(n87), .B2(n187), .A(n84), .ZN(n82) );
  INV_X1 U203 ( .A(n86), .ZN(n84) );
  NOR2_X1 U204 ( .A1(B[3]), .A2(A[3]), .ZN(n80) );
  OR2_X1 U205 ( .A1(B[4]), .A2(A[4]), .ZN(n188) );
  NAND2_X1 U206 ( .A1(B[3]), .A2(A[3]), .ZN(n81) );
  XOR2_X1 U207 ( .A(n16), .B(n91), .Z(SUM[1]) );
  NAND2_X1 U208 ( .A1(n106), .A2(n89), .ZN(n16) );
  INV_X1 U209 ( .A(n88), .ZN(n106) );
  OAI21_X1 U210 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U211 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U212 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  NAND2_X1 U213 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  NAND2_X1 U214 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  XNOR2_X1 U215 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  AOI21_X2 U216 ( .B1(n188), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U217 ( .A1(A[11]), .A2(B[11]), .ZN(n43) );
  XNOR2_X1 U218 ( .A(n1), .B(n189), .ZN(SUM[11]) );
  AND2_X1 U219 ( .A1(n168), .A2(n43), .ZN(n189) );
  XNOR2_X1 U220 ( .A(n10), .B(n65), .ZN(SUM[7]) );
  OAI21_X1 U221 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  AOI21_X1 U222 ( .B1(n65), .B2(n172), .A(n62), .ZN(n60) );
  XNOR2_X1 U223 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U224 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  NAND2_X1 U225 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  NAND2_X1 U226 ( .A1(n104), .A2(n81), .ZN(n14) );
  NAND2_X1 U227 ( .A1(A[12]), .A2(B[12]), .ZN(n40) );
  INV_X1 U228 ( .A(n38), .ZN(n36) );
  AOI21_X1 U229 ( .B1(n23), .B2(n165), .A(n24), .ZN(n22) );
  AOI21_X1 U230 ( .B1(n94), .B2(n38), .A(n31), .ZN(n29) );
  OAI21_X1 U231 ( .B1(n169), .B2(n43), .A(n40), .ZN(n38) );
  NAND2_X1 U232 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  XNOR2_X1 U233 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  OAI21_X1 U234 ( .B1(n50), .B2(n52), .A(n51), .ZN(n49) );
  XNOR2_X1 U235 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  INV_X1 U236 ( .A(n177), .ZN(n97) );
  NOR2_X1 U237 ( .A1(n177), .A2(n50), .ZN(n45) );
  OAI21_X1 U238 ( .B1(n47), .B2(n51), .A(n48), .ZN(n46) );
  INV_X1 U239 ( .A(n174), .ZN(n52) );
  OAI21_X1 U240 ( .B1(n1), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U241 ( .B1(n1), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U242 ( .B1(n180), .B2(n166), .A(n36), .ZN(n34) );
  OAI21_X1 U243 ( .B1(n42), .B2(n180), .A(n167), .ZN(n41) );
  NAND2_X1 U244 ( .A1(n185), .A2(n172), .ZN(n54) );
  AOI21_X1 U245 ( .B1(n185), .B2(n62), .A(n178), .ZN(n55) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_2_DW01_add_5 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n10, n11, n12, n13, n14, n15, n16, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n36,
         n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n57, n59, n60, n62, n64, n65, n66, n68, n70, n71,
         n72, n73, n74, n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89,
         n91, n93, n94, n96, n97, n98, n102, n104, n106, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187;

  CLKBUF_X1 U127 ( .A(A[12]), .Z(n162) );
  CLKBUF_X1 U128 ( .A(B[12]), .Z(n163) );
  OR2_X1 U129 ( .A1(A[8]), .A2(B[8]), .ZN(n184) );
  OR2_X1 U130 ( .A1(n39), .A2(n42), .ZN(n164) );
  BUF_X1 U131 ( .A(n66), .Z(n165) );
  NOR2_X1 U132 ( .A1(B[12]), .A2(A[12]), .ZN(n166) );
  AOI21_X1 U133 ( .B1(n184), .B2(n62), .A(n57), .ZN(n167) );
  INV_X1 U134 ( .A(n96), .ZN(n168) );
  OAI21_X1 U135 ( .B1(n54), .B2(n165), .A(n167), .ZN(n169) );
  BUF_X1 U136 ( .A(n48), .Z(n170) );
  CLKBUF_X1 U137 ( .A(n37), .Z(n171) );
  AND2_X1 U138 ( .A1(n180), .A2(n91), .ZN(SUM[0]) );
  XNOR2_X1 U139 ( .A(n169), .B(n173), .ZN(SUM[9]) );
  NAND2_X1 U140 ( .A1(n98), .A2(n51), .ZN(n173) );
  CLKBUF_X1 U141 ( .A(n38), .Z(n174) );
  XNOR2_X1 U142 ( .A(n179), .B(n175), .ZN(SUM[11]) );
  AND2_X1 U143 ( .A1(n96), .A2(n43), .ZN(n175) );
  CLKBUF_X1 U144 ( .A(n179), .Z(n176) );
  OAI21_X1 U145 ( .B1(n54), .B2(n165), .A(n55), .ZN(n53) );
  INV_X1 U146 ( .A(n50), .ZN(n98) );
  OR2_X1 U147 ( .A1(n163), .A2(n162), .ZN(n177) );
  AOI21_X1 U148 ( .B1(n45), .B2(n53), .A(n46), .ZN(n179) );
  NOR2_X1 U149 ( .A1(B[10]), .A2(A[10]), .ZN(n178) );
  AOI21_X1 U150 ( .B1(n169), .B2(n45), .A(n46), .ZN(n1) );
  OR2_X1 U151 ( .A1(B[7]), .A2(A[7]), .ZN(n185) );
  OR2_X1 U152 ( .A1(B[0]), .A2(A[0]), .ZN(n180) );
  INV_X1 U153 ( .A(n66), .ZN(n65) );
  XNOR2_X1 U154 ( .A(n11), .B(n71), .ZN(SUM[6]) );
  NAND2_X1 U155 ( .A1(n186), .A2(n70), .ZN(n11) );
  INV_X1 U156 ( .A(n42), .ZN(n96) );
  INV_X1 U157 ( .A(n70), .ZN(n68) );
  INV_X1 U158 ( .A(n59), .ZN(n57) );
  NOR2_X1 U159 ( .A1(B[9]), .A2(A[9]), .ZN(n50) );
  XNOR2_X1 U160 ( .A(n60), .B(n181), .ZN(SUM[8]) );
  AND2_X1 U161 ( .A1(n184), .A2(n59), .ZN(n181) );
  XNOR2_X1 U162 ( .A(n49), .B(n7), .ZN(SUM[10]) );
  NAND2_X1 U163 ( .A1(n97), .A2(n170), .ZN(n7) );
  XOR2_X1 U164 ( .A(n12), .B(n74), .Z(SUM[5]) );
  NAND2_X1 U165 ( .A1(n102), .A2(n73), .ZN(n12) );
  INV_X1 U166 ( .A(n72), .ZN(n102) );
  OAI21_X1 U167 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  INV_X1 U168 ( .A(n33), .ZN(n31) );
  NAND2_X1 U169 ( .A1(n93), .A2(n26), .ZN(n3) );
  INV_X1 U170 ( .A(n25), .ZN(n93) );
  NAND2_X1 U171 ( .A1(n177), .A2(n40), .ZN(n5) );
  NAND2_X1 U172 ( .A1(n94), .A2(n33), .ZN(n4) );
  INV_X1 U173 ( .A(n38), .ZN(n36) );
  XNOR2_X1 U174 ( .A(n10), .B(n65), .ZN(SUM[7]) );
  NAND2_X1 U175 ( .A1(n185), .A2(n64), .ZN(n10) );
  XNOR2_X1 U176 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U177 ( .A1(n182), .A2(n19), .ZN(n2) );
  NAND2_X1 U178 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  INV_X1 U179 ( .A(n32), .ZN(n94) );
  NOR2_X1 U180 ( .A1(n32), .A2(n25), .ZN(n23) );
  OR2_X1 U181 ( .A1(B[15]), .A2(A[15]), .ZN(n182) );
  NOR2_X1 U182 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  INV_X1 U183 ( .A(n78), .ZN(n76) );
  XOR2_X1 U184 ( .A(n14), .B(n82), .Z(SUM[3]) );
  NAND2_X1 U185 ( .A1(n104), .A2(n81), .ZN(n14) );
  INV_X1 U186 ( .A(n80), .ZN(n104) );
  NOR2_X1 U187 ( .A1(B[10]), .A2(A[10]), .ZN(n47) );
  NOR2_X1 U188 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  NOR2_X1 U189 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  OAI21_X1 U190 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  OR2_X1 U191 ( .A1(B[2]), .A2(A[2]), .ZN(n183) );
  NAND2_X1 U192 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  NAND2_X1 U193 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  NOR2_X1 U194 ( .A1(B[11]), .A2(A[11]), .ZN(n42) );
  NAND2_X1 U195 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  NAND2_X1 U196 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND2_X1 U197 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U198 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  NAND2_X1 U199 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  OR2_X1 U200 ( .A1(B[6]), .A2(A[6]), .ZN(n186) );
  XNOR2_X1 U201 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  NAND2_X1 U202 ( .A1(n187), .A2(n78), .ZN(n13) );
  NOR2_X1 U203 ( .A1(B[3]), .A2(A[3]), .ZN(n80) );
  AOI21_X1 U204 ( .B1(n87), .B2(n183), .A(n84), .ZN(n82) );
  INV_X1 U205 ( .A(n86), .ZN(n84) );
  NAND2_X1 U206 ( .A1(B[3]), .A2(A[3]), .ZN(n81) );
  NAND2_X1 U207 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  OR2_X1 U208 ( .A1(B[4]), .A2(A[4]), .ZN(n187) );
  XNOR2_X1 U209 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U210 ( .A1(n183), .A2(n86), .ZN(n15) );
  XOR2_X1 U211 ( .A(n16), .B(n91), .Z(SUM[1]) );
  NAND2_X1 U212 ( .A1(n106), .A2(n89), .ZN(n16) );
  INV_X1 U213 ( .A(n88), .ZN(n106) );
  OAI21_X1 U214 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U215 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U216 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  NAND2_X1 U217 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  AOI21_X1 U218 ( .B1(n187), .B2(n79), .A(n76), .ZN(n74) );
  NAND2_X1 U219 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  NOR2_X1 U220 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  NOR2_X1 U221 ( .A1(n39), .A2(n42), .ZN(n37) );
  OAI21_X1 U222 ( .B1(n166), .B2(n43), .A(n40), .ZN(n38) );
  XNOR2_X1 U223 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  AOI21_X1 U224 ( .B1(n186), .B2(n71), .A(n68), .ZN(n66) );
  OAI21_X1 U225 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  AOI21_X1 U226 ( .B1(n65), .B2(n185), .A(n62), .ZN(n60) );
  NAND2_X1 U227 ( .A1(n37), .A2(n94), .ZN(n28) );
  AOI21_X1 U228 ( .B1(n38), .B2(n94), .A(n31), .ZN(n29) );
  NAND2_X1 U229 ( .A1(n171), .A2(n23), .ZN(n21) );
  AOI21_X1 U230 ( .B1(n23), .B2(n174), .A(n24), .ZN(n22) );
  INV_X1 U231 ( .A(n178), .ZN(n97) );
  NOR2_X1 U232 ( .A1(n178), .A2(n50), .ZN(n45) );
  OAI21_X1 U233 ( .B1(n47), .B2(n51), .A(n48), .ZN(n46) );
  NAND2_X1 U234 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  XNOR2_X1 U235 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  OAI21_X1 U236 ( .B1(n52), .B2(n50), .A(n51), .ZN(n49) );
  NAND2_X1 U237 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  XNOR2_X1 U238 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  INV_X1 U239 ( .A(n64), .ZN(n62) );
  INV_X1 U240 ( .A(n53), .ZN(n52) );
  OAI21_X1 U241 ( .B1(n176), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U242 ( .B1(n179), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U243 ( .B1(n1), .B2(n168), .A(n43), .ZN(n41) );
  OAI21_X1 U244 ( .B1(n1), .B2(n164), .A(n36), .ZN(n34) );
  AOI21_X1 U245 ( .B1(n184), .B2(n62), .A(n57), .ZN(n55) );
  NAND2_X1 U246 ( .A1(n184), .A2(n185), .ZN(n54) );
  NAND2_X1 U247 ( .A1(B[8]), .A2(A[8]), .ZN(n59) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_2 ( .in({\in[3][15] , 
        \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , \in[3][10] , 
        \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , \in[3][5] , \in[3][4] , 
        \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , \in[2][15] , 
        \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , \in[2][10] , 
        \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , \in[2][5] , \in[2][4] , 
        \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , \in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \genblk1.inter[1][15] , \genblk1.inter[1][14] ,
         \genblk1.inter[1][13] , \genblk1.inter[1][12] ,
         \genblk1.inter[1][11] , \genblk1.inter[1][10] , \genblk1.inter[1][9] ,
         \genblk1.inter[1][8] , \genblk1.inter[1][7] , \genblk1.inter[1][6] ,
         \genblk1.inter[1][5] , \genblk1.inter[1][4] , \genblk1.inter[1][3] ,
         \genblk1.inter[1][2] , \genblk1.inter[1][1] , \genblk1.inter[1][0] ,
         \genblk1.inter[0][15] , \genblk1.inter[0][14] ,
         \genblk1.inter[0][13] , \genblk1.inter[0][12] ,
         \genblk1.inter[0][11] , \genblk1.inter[0][10] , \genblk1.inter[0][9] ,
         \genblk1.inter[0][8] , \genblk1.inter[0][7] , \genblk1.inter[0][6] ,
         \genblk1.inter[0][5] , \genblk1.inter[0][4] , \genblk1.inter[0][3] ,
         \genblk1.inter[0][2] , \genblk1.inter[0][1] , \genblk1.inter[0][0] ;

  recursive_add_layer_INPUT_SCALE2_WIDTH16_2 \genblk1.next_layer  ( .in({
        \genblk1.inter[1][15] , \genblk1.inter[1][14] , \genblk1.inter[1][13] , 
        \genblk1.inter[1][12] , \genblk1.inter[1][11] , \genblk1.inter[1][10] , 
        \genblk1.inter[1][9] , \genblk1.inter[1][8] , \genblk1.inter[1][7] , 
        \genblk1.inter[1][6] , \genblk1.inter[1][5] , \genblk1.inter[1][4] , 
        \genblk1.inter[1][3] , \genblk1.inter[1][2] , \genblk1.inter[1][1] , 
        \genblk1.inter[1][0] , \genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }), .out(out) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_2_DW01_add_4 add_64_G2 ( .A({
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] }), .B({\in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] }), .CI(1'b0), .SUM({\genblk1.inter[1][15] , \genblk1.inter[1][14] , 
        \genblk1.inter[1][13] , \genblk1.inter[1][12] , \genblk1.inter[1][11] , 
        \genblk1.inter[1][10] , \genblk1.inter[1][9] , \genblk1.inter[1][8] , 
        \genblk1.inter[1][7] , \genblk1.inter[1][6] , \genblk1.inter[1][5] , 
        \genblk1.inter[1][4] , \genblk1.inter[1][3] , \genblk1.inter[1][2] , 
        \genblk1.inter[1][1] , \genblk1.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_2_DW01_add_5 add_64 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM({\genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }) );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_2 ( .a({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , 
        \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , 
        \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , 
        \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , \x[1][7] , 
        \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , 
        \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , 
        \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \multout[3][15] , \multout[3][14] , \multout[3][13] ,
         \multout[3][12] , \multout[3][11] , \multout[3][10] , \multout[3][9] ,
         \multout[3][8] , \multout[3][7] , \multout[3][6] , \multout[3][5] ,
         \multout[3][4] , \multout[3][3] , \multout[3][2] , \multout[3][1] ,
         \multout[3][0] , \multout[2][15] , \multout[2][14] , \multout[2][13] ,
         \multout[2][12] , \multout[2][11] , \multout[2][10] , \multout[2][9] ,
         \multout[2][8] , \multout[2][7] , \multout[2][6] , \multout[2][5] ,
         \multout[2][4] , \multout[2][3] , \multout[2][2] , \multout[2][1] ,
         \multout[2][0] , \multout[1][15] , \multout[1][14] , \multout[1][13] ,
         \multout[1][12] , \multout[1][11] , \multout[1][10] , \multout[1][9] ,
         \multout[1][8] , \multout[1][7] , \multout[1][6] , \multout[1][5] ,
         \multout[1][4] , \multout[1][3] , \multout[1][2] , \multout[1][1] ,
         \multout[1][0] , \multout[0][15] , \multout[0][14] , \multout[0][13] ,
         \multout[0][12] , \multout[0][11] , \multout[0][10] , \multout[0][9] ,
         \multout[0][8] , \multout[0][7] , \multout[0][6] , \multout[0][5] ,
         \multout[0][4] , \multout[0][3] , \multout[0][2] , \multout[0][1] ,
         \multout[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_8 \genblk1[0].mult  ( .ia({\a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({\multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_7 \genblk1[1].mult  ( .ia({\a[1][7] , 
        \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , 
        \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , 
        \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({\multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_6 \genblk1[2].mult  ( .ia({\a[2][7] , 
        \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , \a[2][1] , 
        \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] , 
        \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({\multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_5 \genblk1[3].mult  ( .ia({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_2 add ( .in({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] , \multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] , \multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] , \multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }), .out(y) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n12, n13, n14, n16, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50, n51,
         n52, n53, n56, n58, n61, n62, n63, n64, n65, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n80, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102, n103, n104,
         n105, n108, n109, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n163, n164, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n245, n246, n247, n248, n250, n251, n252,
         n253, n254, n255, n256, n258, n259, n260, n261, n262, n263, n264,
         n265, n273, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n355, n356;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n321), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n195), .B(n188), .CI(n182), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n148), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  XNOR2_X1 U268 ( .A(n133), .B(n303), .ZN(n131) );
  XNOR2_X1 U269 ( .A(n138), .B(n135), .ZN(n303) );
  XOR2_X1 U270 ( .A(b[5]), .B(n261), .Z(n231) );
  CLKBUF_X1 U271 ( .A(n190), .Z(n304) );
  OR2_X1 U272 ( .A1(n143), .A2(n146), .ZN(n305) );
  NAND2_X1 U273 ( .A1(n264), .A2(n307), .ZN(n308) );
  NAND2_X1 U274 ( .A1(n306), .A2(a[2]), .ZN(n309) );
  NAND2_X1 U275 ( .A1(n308), .A2(n309), .ZN(n248) );
  INV_X1 U276 ( .A(n264), .ZN(n306) );
  INV_X1 U277 ( .A(a[2]), .ZN(n307) );
  CLKBUF_X1 U278 ( .A(n89), .Z(n310) );
  CLKBUF_X1 U279 ( .A(n264), .Z(n311) );
  OR2_X2 U280 ( .A1(n312), .A2(n164), .ZN(n253) );
  XNOR2_X1 U281 ( .A(n265), .B(n164), .ZN(n312) );
  INV_X1 U282 ( .A(n164), .ZN(n273) );
  NAND2_X1 U283 ( .A1(n133), .A2(n138), .ZN(n313) );
  NAND2_X1 U284 ( .A1(n133), .A2(n135), .ZN(n314) );
  NAND2_X1 U285 ( .A1(n138), .A2(n135), .ZN(n315) );
  NAND3_X1 U286 ( .A1(n313), .A2(n314), .A3(n315), .ZN(n130) );
  OR2_X1 U287 ( .A1(n229), .A2(n253), .ZN(n316) );
  OR2_X1 U288 ( .A1(n229), .A2(n273), .ZN(n317) );
  NAND2_X1 U289 ( .A1(n316), .A2(n317), .ZN(n163) );
  XNOR2_X1 U290 ( .A(n263), .B(a[6]), .ZN(n318) );
  BUF_X2 U291 ( .A(n256), .Z(n355) );
  CLKBUF_X3 U292 ( .A(n245), .Z(n356) );
  BUF_X1 U293 ( .A(n70), .Z(n319) );
  NOR2_X1 U294 ( .A1(n121), .A2(n124), .ZN(n320) );
  OAI22_X1 U295 ( .A1(n344), .A2(n221), .B1(n220), .B2(n355), .ZN(n321) );
  OR2_X1 U296 ( .A1(n64), .A2(n61), .ZN(n322) );
  NOR2_X1 U297 ( .A1(n334), .A2(n72), .ZN(n67) );
  INV_X1 U298 ( .A(n88), .ZN(n109) );
  BUF_X2 U299 ( .A(n350), .Z(n329) );
  XOR2_X1 U300 ( .A(n190), .B(n197), .Z(n323) );
  XOR2_X1 U301 ( .A(n149), .B(n323), .Z(n147) );
  NAND2_X1 U302 ( .A1(n149), .A2(n304), .ZN(n324) );
  NAND2_X1 U303 ( .A1(n149), .A2(n197), .ZN(n325) );
  NAND2_X1 U304 ( .A1(n190), .A2(n197), .ZN(n326) );
  NAND3_X1 U305 ( .A1(n324), .A2(n325), .A3(n326), .ZN(n146) );
  OAI21_X1 U306 ( .B1(n61), .B2(n65), .A(n62), .ZN(n327) );
  BUF_X1 U307 ( .A(n350), .Z(n328) );
  INV_X1 U308 ( .A(n72), .ZN(n105) );
  OAI21_X1 U309 ( .B1(n320), .B2(n65), .A(n62), .ZN(n2) );
  OR2_X1 U310 ( .A1(n201), .A2(n169), .ZN(n330) );
  XNOR2_X1 U311 ( .A(n264), .B(a[4]), .ZN(n331) );
  CLKBUF_X1 U312 ( .A(n265), .Z(n332) );
  XNOR2_X1 U313 ( .A(n265), .B(a[2]), .ZN(n333) );
  NOR2_X1 U314 ( .A1(n131), .A2(n136), .ZN(n334) );
  NAND2_X1 U315 ( .A1(n246), .A2(n254), .ZN(n335) );
  NOR2_X1 U316 ( .A1(n131), .A2(n136), .ZN(n69) );
  NAND2_X1 U317 ( .A1(n246), .A2(n254), .ZN(n250) );
  XNOR2_X1 U318 ( .A(n264), .B(a[4]), .ZN(n336) );
  INV_X1 U319 ( .A(n260), .ZN(n337) );
  XNOR2_X1 U320 ( .A(n263), .B(a[6]), .ZN(n350) );
  CLKBUF_X1 U321 ( .A(n78), .Z(n338) );
  CLKBUF_X1 U322 ( .A(n262), .Z(n339) );
  CLKBUF_X1 U323 ( .A(n263), .Z(n340) );
  CLKBUF_X1 U324 ( .A(n265), .Z(n341) );
  XNOR2_X1 U325 ( .A(n349), .B(n342), .ZN(product[9]) );
  AND2_X1 U326 ( .A1(n103), .A2(n65), .ZN(n342) );
  BUF_X1 U327 ( .A(n75), .Z(n343) );
  NAND2_X1 U328 ( .A1(n248), .A2(n256), .ZN(n344) );
  NAND2_X1 U329 ( .A1(n248), .A2(n333), .ZN(n345) );
  NAND2_X1 U330 ( .A1(n331), .A2(n247), .ZN(n346) );
  XOR2_X1 U331 ( .A(n347), .B(n90), .Z(product[3]) );
  NAND2_X1 U332 ( .A1(n109), .A2(n310), .ZN(n347) );
  NOR2_X1 U333 ( .A1(n137), .A2(n142), .ZN(n72) );
  NOR2_X1 U334 ( .A1(n121), .A2(n124), .ZN(n61) );
  AOI21_X1 U335 ( .B1(n67), .B2(n343), .A(n68), .ZN(n348) );
  AOI21_X1 U336 ( .B1(n67), .B2(n343), .A(n68), .ZN(n349) );
  INV_X1 U337 ( .A(n30), .ZN(n28) );
  INV_X1 U338 ( .A(n64), .ZN(n103) );
  INV_X1 U339 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U340 ( .A1(n3), .A2(n21), .ZN(n19) );
  AOI21_X1 U341 ( .B1(n2), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U342 ( .B1(n327), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U343 ( .A(n31), .ZN(n29) );
  NAND2_X1 U344 ( .A1(n3), .A2(n39), .ZN(n37) );
  NAND2_X1 U345 ( .A1(n3), .A2(n28), .ZN(n26) );
  NAND2_X1 U346 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U347 ( .A(n41), .ZN(n100) );
  XNOR2_X1 U348 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U349 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U350 ( .A(n34), .ZN(n99) );
  XNOR2_X1 U351 ( .A(n13), .B(n83), .ZN(product[5]) );
  NAND2_X1 U352 ( .A1(n352), .A2(n82), .ZN(n13) );
  NOR2_X1 U353 ( .A1(n64), .A2(n61), .ZN(n3) );
  XNOR2_X1 U354 ( .A(n74), .B(n351), .ZN(product[7]) );
  AND2_X1 U355 ( .A1(n105), .A2(n73), .ZN(n351) );
  XNOR2_X1 U356 ( .A(n56), .B(n7), .ZN(product[11]) );
  INV_X1 U357 ( .A(n2), .ZN(n58) );
  NAND2_X1 U358 ( .A1(n104), .A2(n319), .ZN(n10) );
  OAI21_X1 U359 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  INV_X1 U360 ( .A(n334), .ZN(n104) );
  NAND2_X1 U361 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U362 ( .A(n23), .ZN(n98) );
  AOI21_X1 U363 ( .B1(n352), .B2(n83), .A(n80), .ZN(n78) );
  INV_X1 U364 ( .A(n82), .ZN(n80) );
  AOI21_X1 U365 ( .B1(n353), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U366 ( .A(n94), .ZN(n92) );
  AOI21_X1 U367 ( .B1(n67), .B2(n343), .A(n68), .ZN(n1) );
  AOI21_X1 U368 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U369 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U370 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U371 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U372 ( .A(n320), .ZN(n102) );
  OAI21_X1 U373 ( .B1(n76), .B2(n78), .A(n77), .ZN(n75) );
  NOR2_X1 U374 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U375 ( .A1(n125), .A2(n130), .ZN(n64) );
  NOR2_X1 U376 ( .A1(n50), .A2(n41), .ZN(n39) );
  OAI21_X1 U377 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  NOR2_X1 U378 ( .A1(n41), .A2(n34), .ZN(n32) );
  NAND2_X1 U379 ( .A1(n125), .A2(n130), .ZN(n65) );
  AOI21_X1 U380 ( .B1(n327), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U381 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  INV_X1 U382 ( .A(n51), .ZN(n53) );
  NAND2_X1 U383 ( .A1(n131), .A2(n136), .ZN(n70) );
  INV_X1 U384 ( .A(n50), .ZN(n52) );
  XNOR2_X1 U385 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U386 ( .A1(n353), .A2(n94), .ZN(n16) );
  NAND2_X1 U387 ( .A1(n305), .A2(n77), .ZN(n12) );
  NOR2_X1 U388 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U389 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U390 ( .A1(n187), .A2(n175), .ZN(n134) );
  OAI21_X1 U391 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  NOR2_X1 U392 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U393 ( .A1(n114), .A2(n113), .ZN(n34) );
  INV_X1 U394 ( .A(n112), .ZN(n113) );
  OR2_X1 U395 ( .A1(n147), .A2(n150), .ZN(n352) );
  OAI21_X1 U396 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NOR2_X1 U397 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U398 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U399 ( .A1(n116), .A2(n115), .ZN(n44) );
  INV_X1 U400 ( .A(n97), .ZN(n95) );
  OR2_X1 U401 ( .A1(n200), .A2(n193), .ZN(n353) );
  NOR2_X1 U402 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U403 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U404 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U405 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U406 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U407 ( .A1(n143), .A2(n146), .ZN(n77) );
  AND2_X1 U408 ( .A1(n356), .A2(n161), .ZN(n193) );
  XOR2_X1 U409 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U410 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U411 ( .A(n84), .ZN(n108) );
  OR2_X1 U412 ( .A1(n356), .A2(n259), .ZN(n219) );
  AND2_X1 U413 ( .A1(n356), .A2(n155), .ZN(n177) );
  INV_X1 U414 ( .A(n157), .ZN(n178) );
  AND2_X1 U415 ( .A1(n356), .A2(n158), .ZN(n185) );
  INV_X1 U416 ( .A(n118), .ZN(n119) );
  NOR2_X1 U417 ( .A1(n153), .A2(n168), .ZN(n88) );
  NOR2_X1 U418 ( .A1(n151), .A2(n152), .ZN(n84) );
  INV_X1 U419 ( .A(n163), .ZN(n194) );
  INV_X1 U420 ( .A(n154), .ZN(n170) );
  NAND2_X1 U421 ( .A1(n151), .A2(n152), .ZN(n85) );
  INV_X1 U422 ( .A(n128), .ZN(n129) );
  OR2_X1 U423 ( .A1(n356), .A2(n258), .ZN(n210) );
  AND2_X1 U424 ( .A1(n330), .A2(n97), .ZN(product[1]) );
  XNOR2_X1 U425 ( .A(n263), .B(a[6]), .ZN(n254) );
  OR2_X1 U426 ( .A1(n356), .A2(n260), .ZN(n228) );
  OR2_X1 U427 ( .A1(n356), .A2(n261), .ZN(n237) );
  NAND2_X1 U428 ( .A1(n248), .A2(n256), .ZN(n252) );
  NAND2_X1 U429 ( .A1(n247), .A2(n331), .ZN(n251) );
  AND2_X1 U430 ( .A1(n356), .A2(n164), .ZN(product[0]) );
  INV_X1 U431 ( .A(n160), .ZN(n186) );
  XNOR2_X1 U432 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U433 ( .A(b[7]), .B(n339), .ZN(n202) );
  XNOR2_X1 U434 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U435 ( .A(b[6]), .B(n262), .ZN(n203) );
  XNOR2_X1 U436 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U437 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U438 ( .A(n262), .B(n356), .ZN(n209) );
  INV_X1 U439 ( .A(n262), .ZN(n258) );
  XNOR2_X1 U440 ( .A(b[1]), .B(n262), .ZN(n208) );
  XOR2_X1 U441 ( .A(a[6]), .B(n262), .Z(n246) );
  OAI22_X1 U442 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  OAI22_X1 U443 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  OAI22_X1 U444 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U445 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U446 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U447 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  XNOR2_X1 U448 ( .A(n264), .B(a[4]), .ZN(n255) );
  XNOR2_X1 U449 ( .A(n265), .B(a[2]), .ZN(n256) );
  NAND2_X1 U450 ( .A1(n147), .A2(n150), .ZN(n82) );
  INV_X1 U451 ( .A(n87), .ZN(n86) );
  XNOR2_X1 U452 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U453 ( .A1(n52), .A2(n51), .ZN(n7) );
  NAND2_X1 U454 ( .A1(n3), .A2(n52), .ZN(n46) );
  AOI21_X1 U455 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  NAND2_X1 U456 ( .A1(n52), .A2(n32), .ZN(n30) );
  OAI21_X1 U457 ( .B1(n73), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U458 ( .A(n75), .ZN(n74) );
  XNOR2_X1 U459 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U460 ( .A1(n200), .A2(n193), .ZN(n94) );
  XOR2_X1 U461 ( .A(n12), .B(n338), .Z(product[6]) );
  OAI22_X1 U462 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OAI21_X1 U463 ( .B1(n349), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U464 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  OAI21_X1 U465 ( .B1(n348), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U466 ( .B1(n348), .B2(n322), .A(n58), .ZN(n56) );
  OAI21_X1 U467 ( .B1(n348), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U468 ( .B1(n349), .B2(n26), .A(n27), .ZN(n25) );
  OAI22_X1 U469 ( .A1(n202), .A2(n335), .B1(n202), .B2(n254), .ZN(n154) );
  OAI22_X1 U470 ( .A1(n335), .A2(n206), .B1(n205), .B2(n318), .ZN(n173) );
  OAI22_X1 U471 ( .A1(n335), .A2(n203), .B1(n202), .B2(n318), .ZN(n112) );
  OAI22_X1 U472 ( .A1(n335), .A2(n205), .B1(n204), .B2(n329), .ZN(n172) );
  OAI22_X1 U473 ( .A1(n335), .A2(n204), .B1(n203), .B2(n329), .ZN(n171) );
  OAI22_X1 U474 ( .A1(n335), .A2(n208), .B1(n207), .B2(n318), .ZN(n175) );
  OAI22_X1 U475 ( .A1(n335), .A2(n207), .B1(n206), .B2(n329), .ZN(n174) );
  INV_X1 U476 ( .A(n328), .ZN(n155) );
  XNOR2_X1 U477 ( .A(b[2]), .B(n340), .ZN(n216) );
  OAI22_X1 U478 ( .A1(n250), .A2(n258), .B1(n210), .B2(n318), .ZN(n166) );
  OAI22_X1 U479 ( .A1(n250), .A2(n209), .B1(n208), .B2(n329), .ZN(n176) );
  XNOR2_X1 U480 ( .A(n263), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U481 ( .A(b[3]), .B(n263), .ZN(n215) );
  XNOR2_X1 U482 ( .A(n263), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U483 ( .A(b[4]), .B(n340), .ZN(n214) );
  XNOR2_X1 U484 ( .A(b[7]), .B(n340), .ZN(n211) );
  XNOR2_X1 U485 ( .A(n263), .B(n356), .ZN(n218) );
  XNOR2_X1 U486 ( .A(b[1]), .B(n263), .ZN(n217) );
  INV_X1 U487 ( .A(n263), .ZN(n259) );
  XOR2_X1 U488 ( .A(n263), .B(a[4]), .Z(n247) );
  NAND2_X1 U489 ( .A1(n153), .A2(n168), .ZN(n89) );
  XNOR2_X1 U490 ( .A(b[6]), .B(n265), .ZN(n230) );
  XNOR2_X1 U491 ( .A(b[4]), .B(n341), .ZN(n232) );
  XNOR2_X1 U492 ( .A(n332), .B(n356), .ZN(n236) );
  INV_X1 U493 ( .A(n265), .ZN(n261) );
  XNOR2_X1 U494 ( .A(b[7]), .B(n332), .ZN(n229) );
  XNOR2_X1 U495 ( .A(b[1]), .B(n265), .ZN(n235) );
  XNOR2_X1 U496 ( .A(b[2]), .B(n265), .ZN(n234) );
  XNOR2_X1 U497 ( .A(b[3]), .B(n341), .ZN(n233) );
  NAND2_X1 U498 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U499 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  XNOR2_X1 U500 ( .A(n71), .B(n10), .ZN(product[8]) );
  OAI22_X1 U501 ( .A1(n346), .A2(n217), .B1(n216), .B2(n336), .ZN(n183) );
  OAI22_X1 U502 ( .A1(n346), .A2(n212), .B1(n211), .B2(n255), .ZN(n118) );
  OAI22_X1 U503 ( .A1(n211), .A2(n346), .B1(n211), .B2(n336), .ZN(n157) );
  OAI22_X1 U504 ( .A1(n346), .A2(n213), .B1(n212), .B2(n336), .ZN(n179) );
  OAI22_X1 U505 ( .A1(n346), .A2(n214), .B1(n213), .B2(n255), .ZN(n180) );
  OAI22_X1 U506 ( .A1(n346), .A2(n216), .B1(n215), .B2(n336), .ZN(n182) );
  OAI22_X1 U507 ( .A1(n346), .A2(n215), .B1(n214), .B2(n255), .ZN(n181) );
  INV_X1 U508 ( .A(n255), .ZN(n158) );
  XNOR2_X1 U509 ( .A(b[4]), .B(n264), .ZN(n223) );
  XNOR2_X1 U510 ( .A(n311), .B(b[6]), .ZN(n221) );
  XNOR2_X1 U511 ( .A(b[5]), .B(n337), .ZN(n222) );
  XNOR2_X1 U512 ( .A(b[3]), .B(n264), .ZN(n224) );
  OAI22_X1 U513 ( .A1(n251), .A2(n259), .B1(n219), .B2(n255), .ZN(n167) );
  OAI22_X1 U514 ( .A1(n251), .A2(n218), .B1(n217), .B2(n336), .ZN(n184) );
  XNOR2_X1 U515 ( .A(b[7]), .B(n264), .ZN(n220) );
  XNOR2_X1 U516 ( .A(b[2]), .B(n337), .ZN(n225) );
  INV_X1 U517 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U518 ( .A(n264), .B(n356), .ZN(n227) );
  XNOR2_X1 U519 ( .A(b[1]), .B(n264), .ZN(n226) );
  OAI22_X1 U520 ( .A1(n344), .A2(n221), .B1(n220), .B2(n355), .ZN(n128) );
  OAI22_X1 U521 ( .A1(n220), .A2(n344), .B1(n220), .B2(n333), .ZN(n160) );
  OAI22_X1 U522 ( .A1(n345), .A2(n222), .B1(n221), .B2(n355), .ZN(n187) );
  OAI22_X1 U523 ( .A1(n345), .A2(n223), .B1(n222), .B2(n355), .ZN(n188) );
  OAI22_X1 U524 ( .A1(n344), .A2(n225), .B1(n224), .B2(n355), .ZN(n190) );
  OAI22_X1 U525 ( .A1(n252), .A2(n224), .B1(n223), .B2(n355), .ZN(n189) );
  OAI22_X1 U526 ( .A1(n345), .A2(n226), .B1(n225), .B2(n333), .ZN(n191) );
  OAI22_X1 U527 ( .A1(n344), .A2(n260), .B1(n228), .B2(n333), .ZN(n168) );
  INV_X1 U528 ( .A(n333), .ZN(n161) );
  OAI22_X1 U529 ( .A1(n252), .A2(n227), .B1(n226), .B2(n333), .ZN(n192) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102,
         n103, n105, n108, n109, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n157, n158, n160, n161, n163, n164, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n245, n246, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n258, n259, n260, n261, n262, n263,
         n264, n265, n273, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n341, n342, n343, n344,
         n345, n346;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U136 ( .A(n138), .B(n135), .CI(n133), .CO(n130), .S(n131) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n176), .B(n166), .CO(n140), .S(n141) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n184), .B(n167), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  CLKBUF_X1 U268 ( .A(n263), .Z(n303) );
  AOI21_X1 U269 ( .B1(n322), .B2(n83), .A(n317), .ZN(n304) );
  BUF_X2 U270 ( .A(n262), .Z(n305) );
  BUF_X2 U271 ( .A(n263), .Z(n332) );
  BUF_X2 U272 ( .A(n255), .Z(n344) );
  BUF_X1 U273 ( .A(n264), .Z(n306) );
  BUF_X2 U274 ( .A(n262), .Z(n320) );
  CLKBUF_X1 U275 ( .A(n264), .Z(n307) );
  CLKBUF_X3 U276 ( .A(n245), .Z(n346) );
  CLKBUF_X1 U277 ( .A(n264), .Z(n308) );
  BUF_X2 U278 ( .A(n255), .Z(n345) );
  OR2_X2 U279 ( .A1(n330), .A2(n331), .ZN(n327) );
  BUF_X1 U280 ( .A(n326), .Z(n316) );
  XOR2_X1 U281 ( .A(n148), .B(n183), .Z(n309) );
  XOR2_X1 U282 ( .A(n145), .B(n309), .Z(n143) );
  NAND2_X1 U283 ( .A1(n145), .A2(n148), .ZN(n310) );
  NAND2_X1 U284 ( .A1(n145), .A2(n183), .ZN(n311) );
  NAND2_X1 U285 ( .A1(n148), .A2(n183), .ZN(n312) );
  NAND3_X1 U286 ( .A1(n310), .A2(n311), .A3(n312), .ZN(n142) );
  OR2_X1 U287 ( .A1(n143), .A2(n146), .ZN(n313) );
  XNOR2_X1 U288 ( .A(n303), .B(a[6]), .ZN(n314) );
  XNOR2_X1 U289 ( .A(n263), .B(a[6]), .ZN(n315) );
  XNOR2_X1 U290 ( .A(n263), .B(a[6]), .ZN(n338) );
  AND2_X2 U291 ( .A1(n147), .A2(n150), .ZN(n317) );
  INV_X4 U292 ( .A(n317), .ZN(n82) );
  OAI21_X1 U293 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  INV_X1 U294 ( .A(n260), .ZN(n318) );
  NAND2_X1 U295 ( .A1(n246), .A2(n254), .ZN(n319) );
  NAND2_X1 U296 ( .A1(n246), .A2(n254), .ZN(n250) );
  BUF_X2 U297 ( .A(n256), .Z(n343) );
  FA_X1 U298 ( .A(n138), .B(n135), .CI(n133), .S(n321) );
  OR2_X1 U299 ( .A1(n147), .A2(n150), .ZN(n322) );
  OR2_X1 U300 ( .A1(n201), .A2(n169), .ZN(n323) );
  CLKBUF_X1 U301 ( .A(n304), .Z(n324) );
  NAND2_X1 U302 ( .A1(n248), .A2(n341), .ZN(n325) );
  NAND2_X1 U303 ( .A1(n341), .A2(n248), .ZN(n326) );
  NAND2_X1 U304 ( .A1(n248), .A2(n341), .ZN(n252) );
  CLKBUF_X1 U305 ( .A(n75), .Z(n335) );
  OR2_X1 U306 ( .A1(n330), .A2(n331), .ZN(n251) );
  CLKBUF_X1 U307 ( .A(n265), .Z(n328) );
  CLKBUF_X1 U308 ( .A(n256), .Z(n342) );
  OR2_X1 U309 ( .A1(n321), .A2(n136), .ZN(n329) );
  XOR2_X1 U310 ( .A(n264), .B(a[4]), .Z(n330) );
  XNOR2_X1 U311 ( .A(n263), .B(a[4]), .ZN(n331) );
  CLKBUF_X1 U312 ( .A(n265), .Z(n333) );
  XNOR2_X1 U313 ( .A(n336), .B(n334), .ZN(product[9]) );
  AND2_X1 U314 ( .A1(n103), .A2(n65), .ZN(n334) );
  OAI21_X1 U315 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  XNOR2_X1 U316 ( .A(n13), .B(n83), .ZN(product[5]) );
  XNOR2_X1 U317 ( .A(n56), .B(n7), .ZN(product[11]) );
  AOI21_X1 U318 ( .B1(n67), .B2(n335), .A(n68), .ZN(n336) );
  AOI21_X1 U319 ( .B1(n67), .B2(n335), .A(n68), .ZN(n337) );
  AOI21_X1 U320 ( .B1(n67), .B2(n335), .A(n68), .ZN(n1) );
  XNOR2_X1 U321 ( .A(n263), .B(a[6]), .ZN(n254) );
  NOR2_X1 U322 ( .A1(n121), .A2(n124), .ZN(n61) );
  INV_X1 U323 ( .A(n30), .ZN(n28) );
  INV_X1 U324 ( .A(n64), .ZN(n103) );
  INV_X1 U325 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U326 ( .A1(n3), .A2(n21), .ZN(n19) );
  AOI21_X1 U327 ( .B1(n2), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U328 ( .B1(n2), .B2(n28), .A(n29), .ZN(n27) );
  INV_X1 U329 ( .A(n31), .ZN(n29) );
  NAND2_X1 U330 ( .A1(n3), .A2(n39), .ZN(n37) );
  NAND2_X1 U331 ( .A1(n3), .A2(n28), .ZN(n26) );
  INV_X1 U332 ( .A(n3), .ZN(n57) );
  XNOR2_X1 U333 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U334 ( .A1(n339), .A2(n94), .ZN(n16) );
  NOR2_X1 U335 ( .A1(n64), .A2(n61), .ZN(n3) );
  XNOR2_X1 U336 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U337 ( .A1(n100), .A2(n44), .ZN(n6) );
  INV_X1 U338 ( .A(n41), .ZN(n100) );
  NAND2_X1 U339 ( .A1(n105), .A2(n73), .ZN(n11) );
  INV_X1 U340 ( .A(n72), .ZN(n105) );
  INV_X1 U341 ( .A(n2), .ZN(n58) );
  XNOR2_X1 U342 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U343 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U344 ( .A(n34), .ZN(n99) );
  NAND2_X1 U345 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U346 ( .A(n23), .ZN(n98) );
  AOI21_X1 U347 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U348 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U349 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U350 ( .A1(n102), .A2(n62), .ZN(n8) );
  INV_X1 U351 ( .A(n61), .ZN(n102) );
  NOR2_X1 U352 ( .A1(n30), .A2(n23), .ZN(n21) );
  NOR2_X1 U353 ( .A1(n125), .A2(n130), .ZN(n64) );
  NOR2_X1 U354 ( .A1(n50), .A2(n41), .ZN(n39) );
  AOI21_X1 U355 ( .B1(n339), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U356 ( .A(n94), .ZN(n92) );
  XNOR2_X1 U357 ( .A(n71), .B(n10), .ZN(product[8]) );
  NAND2_X1 U358 ( .A1(n329), .A2(n70), .ZN(n10) );
  OAI21_X1 U359 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  NOR2_X1 U360 ( .A1(n131), .A2(n136), .ZN(n69) );
  NOR2_X1 U361 ( .A1(n41), .A2(n34), .ZN(n32) );
  NAND2_X1 U362 ( .A1(n125), .A2(n130), .ZN(n65) );
  AOI21_X1 U363 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U364 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  INV_X1 U365 ( .A(n51), .ZN(n53) );
  NAND2_X1 U366 ( .A1(n321), .A2(n136), .ZN(n70) );
  INV_X1 U367 ( .A(n50), .ZN(n52) );
  NAND2_X1 U368 ( .A1(n322), .A2(n82), .ZN(n13) );
  NAND2_X1 U369 ( .A1(n313), .A2(n77), .ZN(n12) );
  XOR2_X1 U370 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U371 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U372 ( .A(n84), .ZN(n108) );
  NOR2_X1 U373 ( .A1(n116), .A2(n115), .ZN(n41) );
  XNOR2_X1 U374 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U375 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U376 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U377 ( .A1(n114), .A2(n113), .ZN(n34) );
  XOR2_X1 U378 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U379 ( .A(n88), .ZN(n109) );
  INV_X1 U380 ( .A(n112), .ZN(n113) );
  NOR2_X1 U381 ( .A1(n117), .A2(n120), .ZN(n50) );
  NAND2_X1 U382 ( .A1(n170), .A2(n112), .ZN(n24) );
  NAND2_X1 U383 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U384 ( .A1(n137), .A2(n142), .ZN(n72) );
  INV_X1 U385 ( .A(n97), .ZN(n95) );
  OR2_X1 U386 ( .A1(n200), .A2(n193), .ZN(n339) );
  NOR2_X1 U387 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U388 ( .A1(n121), .A2(n124), .ZN(n62) );
  NAND2_X1 U389 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U390 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U391 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U392 ( .A1(n143), .A2(n146), .ZN(n77) );
  AND2_X1 U393 ( .A1(n346), .A2(n161), .ZN(n193) );
  OAI22_X1 U394 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  AND2_X1 U395 ( .A1(n346), .A2(n158), .ZN(n185) );
  INV_X1 U396 ( .A(n118), .ZN(n119) );
  OR2_X1 U397 ( .A1(n346), .A2(n259), .ZN(n219) );
  OAI22_X1 U398 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  NOR2_X1 U399 ( .A1(n151), .A2(n152), .ZN(n84) );
  INV_X1 U400 ( .A(n128), .ZN(n129) );
  INV_X1 U401 ( .A(n163), .ZN(n194) );
  OAI22_X1 U402 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  OAI22_X1 U403 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  AND2_X1 U404 ( .A1(n346), .A2(n155), .ZN(n177) );
  OAI22_X1 U405 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  NOR2_X1 U406 ( .A1(n153), .A2(n168), .ZN(n88) );
  INV_X1 U407 ( .A(n154), .ZN(n170) );
  NAND2_X1 U408 ( .A1(n151), .A2(n152), .ZN(n85) );
  OR2_X1 U409 ( .A1(n346), .A2(n258), .ZN(n210) );
  INV_X1 U410 ( .A(n157), .ZN(n178) );
  AND2_X1 U411 ( .A1(n323), .A2(n97), .ZN(product[1]) );
  OR2_X1 U412 ( .A1(n346), .A2(n260), .ZN(n228) );
  OAI22_X1 U413 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U414 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OAI22_X1 U415 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OR2_X1 U416 ( .A1(n346), .A2(n261), .ZN(n237) );
  XNOR2_X1 U417 ( .A(b[7]), .B(n305), .ZN(n202) );
  XNOR2_X1 U418 ( .A(b[4]), .B(n320), .ZN(n205) );
  XNOR2_X1 U419 ( .A(b[3]), .B(n320), .ZN(n206) );
  XNOR2_X1 U420 ( .A(b[5]), .B(n305), .ZN(n204) );
  XNOR2_X1 U421 ( .A(b[6]), .B(n320), .ZN(n203) );
  XOR2_X1 U422 ( .A(n262), .B(a[6]), .Z(n246) );
  XNOR2_X1 U423 ( .A(n305), .B(n346), .ZN(n209) );
  INV_X1 U424 ( .A(n262), .ZN(n258) );
  AND2_X1 U425 ( .A1(n346), .A2(n164), .ZN(product[0]) );
  NAND2_X1 U426 ( .A1(n109), .A2(n89), .ZN(n15) );
  OAI21_X1 U427 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  INV_X1 U428 ( .A(n160), .ZN(n186) );
  NAND2_X2 U429 ( .A1(n249), .A2(n273), .ZN(n253) );
  BUF_X1 U430 ( .A(n256), .Z(n341) );
  XNOR2_X1 U431 ( .A(n265), .B(a[2]), .ZN(n256) );
  NAND2_X1 U432 ( .A1(n200), .A2(n193), .ZN(n94) );
  OAI22_X1 U433 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OAI21_X1 U434 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  NOR2_X1 U435 ( .A1(n69), .A2(n72), .ZN(n67) );
  XNOR2_X1 U436 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U437 ( .A1(n52), .A2(n51), .ZN(n7) );
  AOI21_X1 U438 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  NAND2_X1 U439 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U440 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U441 ( .A1(n153), .A2(n168), .ZN(n89) );
  INV_X1 U442 ( .A(n87), .ZN(n86) );
  XNOR2_X1 U443 ( .A(b[2]), .B(n305), .ZN(n207) );
  OAI21_X1 U444 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  XOR2_X1 U445 ( .A(n74), .B(n11), .Z(product[7]) );
  XNOR2_X1 U446 ( .A(n320), .B(b[1]), .ZN(n208) );
  XNOR2_X1 U447 ( .A(b[5]), .B(n318), .ZN(n222) );
  XNOR2_X1 U448 ( .A(b[3]), .B(n308), .ZN(n224) );
  XNOR2_X1 U449 ( .A(b[2]), .B(n307), .ZN(n225) );
  INV_X1 U450 ( .A(n264), .ZN(n260) );
  XNOR2_X1 U451 ( .A(b[6]), .B(n306), .ZN(n221) );
  XNOR2_X1 U452 ( .A(b[4]), .B(n307), .ZN(n223) );
  XNOR2_X1 U453 ( .A(b[7]), .B(n306), .ZN(n220) );
  XNOR2_X1 U454 ( .A(n306), .B(n346), .ZN(n227) );
  XNOR2_X1 U455 ( .A(b[1]), .B(n264), .ZN(n226) );
  XOR2_X1 U456 ( .A(n264), .B(a[2]), .Z(n248) );
  XNOR2_X1 U457 ( .A(n264), .B(a[4]), .ZN(n255) );
  XNOR2_X1 U458 ( .A(n263), .B(n346), .ZN(n218) );
  XNOR2_X1 U459 ( .A(b[1]), .B(n263), .ZN(n217) );
  XNOR2_X1 U460 ( .A(b[2]), .B(n332), .ZN(n216) );
  XNOR2_X1 U461 ( .A(b[3]), .B(n332), .ZN(n215) );
  XNOR2_X1 U462 ( .A(b[4]), .B(n332), .ZN(n214) );
  XNOR2_X1 U463 ( .A(b[5]), .B(n303), .ZN(n213) );
  XNOR2_X1 U464 ( .A(b[6]), .B(n303), .ZN(n212) );
  XNOR2_X1 U465 ( .A(b[7]), .B(n332), .ZN(n211) );
  INV_X1 U466 ( .A(n263), .ZN(n259) );
  AOI21_X1 U467 ( .B1(n322), .B2(n83), .A(n317), .ZN(n78) );
  OAI21_X1 U468 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  XOR2_X1 U469 ( .A(n12), .B(n324), .Z(product[6]) );
  INV_X1 U470 ( .A(n75), .ZN(n74) );
  NAND2_X1 U471 ( .A1(n201), .A2(n169), .ZN(n97) );
  XNOR2_X1 U472 ( .A(b[5]), .B(n333), .ZN(n231) );
  XNOR2_X1 U473 ( .A(b[6]), .B(n333), .ZN(n230) );
  XNOR2_X1 U474 ( .A(b[4]), .B(n333), .ZN(n232) );
  XNOR2_X1 U475 ( .A(b[7]), .B(n328), .ZN(n229) );
  XNOR2_X1 U476 ( .A(n333), .B(n346), .ZN(n236) );
  XNOR2_X1 U477 ( .A(b[3]), .B(n328), .ZN(n233) );
  XNOR2_X1 U478 ( .A(b[2]), .B(n333), .ZN(n234) );
  XNOR2_X1 U479 ( .A(b[1]), .B(n328), .ZN(n235) );
  INV_X1 U480 ( .A(n265), .ZN(n261) );
  XOR2_X1 U481 ( .A(n265), .B(n164), .Z(n249) );
  OAI21_X1 U482 ( .B1(n336), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U483 ( .B1(n336), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U484 ( .B1(n337), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U485 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  OAI21_X1 U486 ( .B1(n337), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U487 ( .B1(n337), .B2(n46), .A(n47), .ZN(n45) );
  OAI22_X1 U488 ( .A1(n202), .A2(n319), .B1(n202), .B2(n314), .ZN(n154) );
  OAI22_X1 U489 ( .A1(n319), .A2(n206), .B1(n205), .B2(n315), .ZN(n173) );
  OAI22_X1 U490 ( .A1(n319), .A2(n203), .B1(n202), .B2(n315), .ZN(n112) );
  OAI22_X1 U491 ( .A1(n319), .A2(n205), .B1(n204), .B2(n314), .ZN(n172) );
  OAI22_X1 U492 ( .A1(n319), .A2(n204), .B1(n203), .B2(n314), .ZN(n171) );
  OAI22_X1 U493 ( .A1(n319), .A2(n208), .B1(n207), .B2(n315), .ZN(n175) );
  OAI22_X1 U494 ( .A1(n319), .A2(n207), .B1(n206), .B2(n314), .ZN(n174) );
  INV_X1 U495 ( .A(n315), .ZN(n155) );
  OAI22_X1 U496 ( .A1(n250), .A2(n258), .B1(n210), .B2(n338), .ZN(n166) );
  OAI22_X1 U497 ( .A1(n250), .A2(n209), .B1(n208), .B2(n338), .ZN(n176) );
  OAI22_X1 U498 ( .A1(n327), .A2(n217), .B1(n216), .B2(n344), .ZN(n183) );
  OAI22_X1 U499 ( .A1(n327), .A2(n212), .B1(n211), .B2(n345), .ZN(n118) );
  OAI22_X1 U500 ( .A1(n211), .A2(n327), .B1(n211), .B2(n345), .ZN(n157) );
  OAI22_X1 U501 ( .A1(n327), .A2(n213), .B1(n212), .B2(n344), .ZN(n179) );
  OAI22_X1 U502 ( .A1(n327), .A2(n214), .B1(n213), .B2(n344), .ZN(n180) );
  OAI22_X1 U503 ( .A1(n327), .A2(n216), .B1(n215), .B2(n345), .ZN(n182) );
  OAI22_X1 U504 ( .A1(n327), .A2(n215), .B1(n214), .B2(n344), .ZN(n181) );
  INV_X1 U505 ( .A(n345), .ZN(n158) );
  OAI22_X1 U506 ( .A1(n251), .A2(n259), .B1(n219), .B2(n345), .ZN(n167) );
  OAI22_X1 U507 ( .A1(n251), .A2(n218), .B1(n217), .B2(n344), .ZN(n184) );
  OAI22_X1 U508 ( .A1(n326), .A2(n221), .B1(n220), .B2(n343), .ZN(n128) );
  OAI22_X1 U509 ( .A1(n220), .A2(n325), .B1(n220), .B2(n343), .ZN(n160) );
  OAI22_X1 U510 ( .A1(n325), .A2(n222), .B1(n221), .B2(n343), .ZN(n187) );
  OAI22_X1 U511 ( .A1(n316), .A2(n224), .B1(n223), .B2(n343), .ZN(n189) );
  OAI22_X1 U512 ( .A1(n325), .A2(n225), .B1(n224), .B2(n342), .ZN(n190) );
  OAI22_X1 U513 ( .A1(n326), .A2(n223), .B1(n222), .B2(n343), .ZN(n188) );
  OAI22_X1 U514 ( .A1(n316), .A2(n260), .B1(n228), .B2(n343), .ZN(n168) );
  OAI22_X1 U515 ( .A1(n325), .A2(n226), .B1(n225), .B2(n342), .ZN(n191) );
  OAI22_X1 U516 ( .A1(n252), .A2(n227), .B1(n226), .B2(n343), .ZN(n192) );
  INV_X1 U517 ( .A(n342), .ZN(n161) );
  INV_X2 U518 ( .A(n164), .ZN(n273) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n50, n51, n52, n53, n56, n58, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n103, n104,
         n108, n109, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n149, n150, n151, n152, n153, n154,
         n155, n157, n160, n161, n163, n164, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n245, n248, n250, n251, n252, n253, n254, n256, n258, n259,
         n260, n261, n262, n263, n264, n265, n273, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n346, n347, n348, n349, n350, n351;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U136 ( .A(n138), .B(n135), .CI(n133), .CO(n130), .S(n131) );
  FA_X1 U137 ( .A(n194), .B(n181), .CI(n140), .CO(n132), .S(n133) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U143 ( .A(n321), .B(n183), .CI(n145), .CO(n142), .S(n143) );
  FA_X1 U144 ( .A(n177), .B(n189), .CI(n196), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n192), .B(n199), .CO(n152), .S(n153) );
  CLKBUF_X3 U268 ( .A(n263), .Z(n350) );
  BUF_X1 U269 ( .A(n348), .Z(n303) );
  CLKBUF_X1 U270 ( .A(n254), .Z(n348) );
  CLKBUF_X1 U271 ( .A(n77), .Z(n304) );
  CLKBUF_X2 U272 ( .A(n262), .Z(n326) );
  OR2_X2 U273 ( .A1(n336), .A2(n337), .ZN(n317) );
  CLKBUF_X1 U274 ( .A(n263), .Z(n305) );
  INV_X1 U275 ( .A(n342), .ZN(n306) );
  OR2_X1 U276 ( .A1(n137), .A2(n142), .ZN(n307) );
  NOR2_X1 U277 ( .A1(n69), .A2(n72), .ZN(n308) );
  BUF_X1 U278 ( .A(n83), .Z(n309) );
  BUF_X2 U279 ( .A(n264), .Z(n310) );
  BUF_X1 U280 ( .A(n262), .Z(n325) );
  OAI21_X1 U281 ( .B1(n61), .B2(n65), .A(n62), .ZN(n311) );
  OR2_X2 U282 ( .A1(n150), .A2(n147), .ZN(n343) );
  NOR2_X1 U283 ( .A1(n131), .A2(n136), .ZN(n312) );
  NOR2_X1 U284 ( .A1(n131), .A2(n136), .ZN(n69) );
  CLKBUF_X1 U285 ( .A(n264), .Z(n313) );
  CLKBUF_X1 U286 ( .A(n264), .Z(n314) );
  OAI21_X1 U287 ( .B1(n312), .B2(n73), .A(n70), .ZN(n315) );
  CLKBUF_X1 U288 ( .A(n265), .Z(n316) );
  OR2_X1 U289 ( .A1(n336), .A2(n337), .ZN(n251) );
  OAI22_X1 U290 ( .A1(n317), .A2(n218), .B1(n217), .B2(n342), .ZN(n318) );
  AOI21_X1 U291 ( .B1(n308), .B2(n339), .A(n315), .ZN(n319) );
  CLKBUF_X1 U292 ( .A(n264), .Z(n320) );
  XNOR2_X2 U293 ( .A(n264), .B(a[4]), .ZN(n342) );
  OAI21_X1 U294 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  AND2_X1 U295 ( .A1(n167), .A2(n318), .ZN(n321) );
  OR2_X1 U296 ( .A1(n201), .A2(n169), .ZN(n322) );
  AND2_X1 U297 ( .A1(n147), .A2(n150), .ZN(n323) );
  AOI21_X1 U298 ( .B1(n343), .B2(n83), .A(n323), .ZN(n324) );
  XOR2_X1 U299 ( .A(a[6]), .B(n325), .Z(n327) );
  INV_X1 U300 ( .A(n265), .ZN(n328) );
  INV_X2 U301 ( .A(n328), .ZN(n329) );
  AOI21_X1 U302 ( .B1(n343), .B2(n83), .A(n323), .ZN(n78) );
  BUF_X1 U303 ( .A(n340), .Z(n330) );
  OR2_X1 U304 ( .A1(n143), .A2(n146), .ZN(n331) );
  OR2_X1 U305 ( .A1(n121), .A2(n124), .ZN(n332) );
  OR2_X1 U306 ( .A1(n64), .A2(n61), .ZN(n333) );
  XOR2_X1 U307 ( .A(n167), .B(n184), .Z(n149) );
  OR2_X2 U308 ( .A1(n334), .A2(n164), .ZN(n253) );
  XNOR2_X1 U309 ( .A(n265), .B(n164), .ZN(n334) );
  INV_X1 U310 ( .A(n164), .ZN(n273) );
  BUF_X1 U311 ( .A(n256), .Z(n346) );
  CLKBUF_X3 U312 ( .A(n256), .Z(n347) );
  AOI21_X1 U313 ( .B1(n67), .B2(n339), .A(n68), .ZN(n335) );
  XOR2_X1 U314 ( .A(n264), .B(a[4]), .Z(n336) );
  XNOR2_X1 U315 ( .A(n263), .B(a[4]), .ZN(n337) );
  XNOR2_X1 U316 ( .A(n1), .B(n338), .ZN(product[9]) );
  AND2_X1 U317 ( .A1(n103), .A2(n65), .ZN(n338) );
  XNOR2_X1 U318 ( .A(n13), .B(n309), .ZN(product[5]) );
  OAI21_X1 U319 ( .B1(n324), .B2(n76), .A(n77), .ZN(n339) );
  NAND2_X1 U320 ( .A1(n248), .A2(n346), .ZN(n340) );
  AOI21_X1 U321 ( .B1(n308), .B2(n339), .A(n315), .ZN(n1) );
  NAND2_X1 U322 ( .A1(n254), .A2(n327), .ZN(n341) );
  NOR2_X1 U323 ( .A1(n64), .A2(n61), .ZN(n3) );
  BUF_X2 U324 ( .A(n245), .Z(n351) );
  NOR2_X1 U325 ( .A1(n151), .A2(n152), .ZN(n84) );
  NAND2_X1 U326 ( .A1(n327), .A2(n254), .ZN(n250) );
  INV_X1 U327 ( .A(n30), .ZN(n28) );
  INV_X1 U328 ( .A(n64), .ZN(n103) );
  INV_X1 U329 ( .A(n31), .ZN(n29) );
  INV_X1 U330 ( .A(n18), .ZN(product[15]) );
  NAND2_X1 U331 ( .A1(n3), .A2(n21), .ZN(n19) );
  NAND2_X1 U332 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U333 ( .A1(n3), .A2(n52), .ZN(n46) );
  NAND2_X1 U334 ( .A1(n3), .A2(n39), .ZN(n37) );
  NAND2_X1 U335 ( .A1(n3), .A2(n28), .ZN(n26) );
  XNOR2_X1 U336 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U337 ( .A1(n99), .A2(n35), .ZN(n5) );
  INV_X1 U338 ( .A(n34), .ZN(n99) );
  XNOR2_X1 U339 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U340 ( .A1(n344), .A2(n94), .ZN(n16) );
  NAND2_X1 U341 ( .A1(n343), .A2(n82), .ZN(n13) );
  NAND2_X1 U342 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U343 ( .A(n23), .ZN(n98) );
  NAND2_X1 U344 ( .A1(n307), .A2(n73), .ZN(n11) );
  XNOR2_X1 U345 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U346 ( .A1(n52), .A2(n51), .ZN(n7) );
  XNOR2_X1 U347 ( .A(n63), .B(n8), .ZN(product[10]) );
  NAND2_X1 U348 ( .A1(n332), .A2(n62), .ZN(n8) );
  NAND2_X1 U349 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U350 ( .A(n69), .ZN(n104) );
  INV_X1 U351 ( .A(n50), .ZN(n52) );
  AOI21_X1 U352 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U353 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U354 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U355 ( .A1(n100), .A2(n44), .ZN(n6) );
  OAI21_X1 U356 ( .B1(n76), .B2(n78), .A(n77), .ZN(n75) );
  NOR2_X1 U357 ( .A1(n125), .A2(n130), .ZN(n64) );
  AOI21_X1 U358 ( .B1(n344), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U359 ( .A(n94), .ZN(n92) );
  NOR2_X1 U360 ( .A1(n30), .A2(n23), .ZN(n21) );
  NAND2_X1 U361 ( .A1(n125), .A2(n130), .ZN(n65) );
  OAI21_X1 U362 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U363 ( .A(n51), .ZN(n53) );
  NAND2_X1 U364 ( .A1(n131), .A2(n136), .ZN(n70) );
  XOR2_X1 U365 ( .A(n12), .B(n324), .Z(product[6]) );
  NAND2_X1 U366 ( .A1(n331), .A2(n304), .ZN(n12) );
  XOR2_X1 U367 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U368 ( .A(n88), .ZN(n109) );
  XNOR2_X1 U369 ( .A(n187), .B(n175), .ZN(n135) );
  OR2_X1 U370 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U371 ( .A1(n170), .A2(n112), .ZN(n23) );
  INV_X1 U372 ( .A(n112), .ZN(n113) );
  NOR2_X1 U373 ( .A1(n121), .A2(n124), .ZN(n61) );
  NOR2_X1 U374 ( .A1(n114), .A2(n113), .ZN(n34) );
  OAI21_X1 U375 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  NAND2_X1 U376 ( .A1(n170), .A2(n112), .ZN(n24) );
  NOR2_X1 U377 ( .A1(n116), .A2(n115), .ZN(n41) );
  NOR2_X1 U378 ( .A1(n137), .A2(n142), .ZN(n72) );
  INV_X1 U379 ( .A(n97), .ZN(n95) );
  OR2_X1 U380 ( .A1(n200), .A2(n193), .ZN(n344) );
  NOR2_X1 U381 ( .A1(n143), .A2(n146), .ZN(n76) );
  NAND2_X1 U382 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U383 ( .A1(n117), .A2(n120), .ZN(n50) );
  INV_X1 U384 ( .A(n87), .ZN(n86) );
  NAND2_X1 U385 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U386 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U387 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U388 ( .A1(n143), .A2(n146), .ZN(n77) );
  NAND2_X1 U389 ( .A1(n121), .A2(n124), .ZN(n62) );
  AND2_X1 U390 ( .A1(n351), .A2(n161), .ZN(n193) );
  XOR2_X1 U391 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U392 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U393 ( .A(n84), .ZN(n108) );
  OR2_X1 U394 ( .A1(n351), .A2(n259), .ZN(n219) );
  INV_X1 U395 ( .A(n157), .ZN(n178) );
  INV_X1 U396 ( .A(n118), .ZN(n119) );
  AND2_X1 U397 ( .A1(n306), .A2(n351), .ZN(n185) );
  OAI22_X1 U398 ( .A1(n253), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U399 ( .A1(n253), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  AND2_X1 U400 ( .A1(n351), .A2(n155), .ZN(n177) );
  OAI22_X1 U401 ( .A1(n253), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U402 ( .A1(n253), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  NOR2_X1 U403 ( .A1(n153), .A2(n168), .ZN(n88) );
  NAND2_X1 U404 ( .A1(n151), .A2(n152), .ZN(n85) );
  INV_X1 U405 ( .A(n154), .ZN(n170) );
  INV_X1 U406 ( .A(n128), .ZN(n129) );
  OR2_X1 U407 ( .A1(n351), .A2(n258), .ZN(n210) );
  AND2_X1 U408 ( .A1(n322), .A2(n97), .ZN(product[1]) );
  INV_X1 U409 ( .A(n163), .ZN(n194) );
  OAI22_X1 U410 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  OR2_X1 U411 ( .A1(n351), .A2(n260), .ZN(n228) );
  OAI22_X1 U412 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U413 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OAI22_X1 U414 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  OR2_X1 U415 ( .A1(n351), .A2(n261), .ZN(n237) );
  NAND2_X1 U416 ( .A1(n248), .A2(n346), .ZN(n252) );
  AND2_X1 U417 ( .A1(n351), .A2(n164), .ZN(product[0]) );
  XNOR2_X1 U418 ( .A(b[4]), .B(n326), .ZN(n205) );
  XNOR2_X1 U419 ( .A(b[7]), .B(n326), .ZN(n202) );
  XNOR2_X1 U420 ( .A(b[6]), .B(n326), .ZN(n203) );
  XNOR2_X1 U421 ( .A(b[5]), .B(n326), .ZN(n204) );
  XNOR2_X1 U422 ( .A(b[2]), .B(n326), .ZN(n207) );
  XNOR2_X1 U423 ( .A(b[3]), .B(n326), .ZN(n206) );
  XNOR2_X1 U424 ( .A(n326), .B(n351), .ZN(n209) );
  INV_X1 U425 ( .A(n325), .ZN(n258) );
  XNOR2_X1 U426 ( .A(b[1]), .B(n326), .ZN(n208) );
  AOI21_X1 U427 ( .B1(n311), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U428 ( .B1(n311), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U429 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U430 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  INV_X1 U431 ( .A(n311), .ZN(n58) );
  INV_X1 U432 ( .A(n160), .ZN(n186) );
  XNOR2_X1 U433 ( .A(n265), .B(a[2]), .ZN(n256) );
  INV_X1 U434 ( .A(n41), .ZN(n100) );
  OAI21_X1 U435 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  NOR2_X1 U436 ( .A1(n50), .A2(n41), .ZN(n39) );
  NOR2_X1 U437 ( .A1(n41), .A2(n34), .ZN(n32) );
  OAI21_X1 U438 ( .B1(n312), .B2(n73), .A(n70), .ZN(n68) );
  NOR2_X1 U439 ( .A1(n69), .A2(n72), .ZN(n67) );
  BUF_X2 U440 ( .A(n254), .Z(n349) );
  XNOR2_X1 U441 ( .A(n263), .B(a[6]), .ZN(n254) );
  XNOR2_X1 U442 ( .A(n25), .B(n4), .ZN(product[14]) );
  XNOR2_X1 U443 ( .A(n71), .B(n10), .ZN(product[8]) );
  NAND2_X1 U444 ( .A1(n109), .A2(n89), .ZN(n15) );
  OAI21_X1 U445 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  XOR2_X1 U446 ( .A(n74), .B(n11), .Z(product[7]) );
  OAI21_X1 U447 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  NAND2_X1 U448 ( .A1(n147), .A2(n150), .ZN(n82) );
  NAND2_X1 U449 ( .A1(n200), .A2(n193), .ZN(n94) );
  INV_X1 U450 ( .A(n75), .ZN(n74) );
  OAI22_X1 U451 ( .A1(n253), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OAI22_X1 U452 ( .A1(n202), .A2(n341), .B1(n202), .B2(n303), .ZN(n154) );
  OAI22_X1 U453 ( .A1(n341), .A2(n203), .B1(n202), .B2(n349), .ZN(n112) );
  OAI22_X1 U454 ( .A1(n341), .A2(n206), .B1(n205), .B2(n349), .ZN(n173) );
  OAI22_X1 U455 ( .A1(n341), .A2(n205), .B1(n204), .B2(n303), .ZN(n172) );
  OAI22_X1 U456 ( .A1(n341), .A2(n204), .B1(n203), .B2(n303), .ZN(n171) );
  OAI22_X1 U457 ( .A1(n341), .A2(n208), .B1(n207), .B2(n349), .ZN(n175) );
  OAI22_X1 U458 ( .A1(n341), .A2(n207), .B1(n206), .B2(n303), .ZN(n174) );
  OAI22_X1 U459 ( .A1(n250), .A2(n258), .B1(n210), .B2(n349), .ZN(n166) );
  OAI22_X1 U460 ( .A1(n250), .A2(n209), .B1(n208), .B2(n348), .ZN(n176) );
  XNOR2_X1 U461 ( .A(b[2]), .B(n350), .ZN(n216) );
  XNOR2_X1 U462 ( .A(b[3]), .B(n350), .ZN(n215) );
  INV_X1 U463 ( .A(n349), .ZN(n155) );
  XNOR2_X1 U464 ( .A(b[7]), .B(n350), .ZN(n211) );
  XNOR2_X1 U465 ( .A(b[4]), .B(n350), .ZN(n214) );
  XNOR2_X1 U466 ( .A(b[5]), .B(n350), .ZN(n213) );
  XNOR2_X1 U467 ( .A(b[6]), .B(n350), .ZN(n212) );
  XNOR2_X1 U468 ( .A(n350), .B(n351), .ZN(n218) );
  INV_X1 U469 ( .A(n305), .ZN(n259) );
  XNOR2_X1 U470 ( .A(b[1]), .B(n350), .ZN(n217) );
  OAI22_X1 U471 ( .A1(n317), .A2(n217), .B1(n216), .B2(n342), .ZN(n183) );
  OAI22_X1 U472 ( .A1(n317), .A2(n212), .B1(n211), .B2(n342), .ZN(n118) );
  OAI22_X1 U473 ( .A1(n211), .A2(n317), .B1(n211), .B2(n342), .ZN(n157) );
  OAI22_X1 U474 ( .A1(n317), .A2(n216), .B1(n215), .B2(n342), .ZN(n182) );
  OAI22_X1 U475 ( .A1(n317), .A2(n214), .B1(n213), .B2(n342), .ZN(n180) );
  OAI22_X1 U476 ( .A1(n317), .A2(n213), .B1(n212), .B2(n342), .ZN(n179) );
  OAI22_X1 U477 ( .A1(n251), .A2(n215), .B1(n214), .B2(n342), .ZN(n181) );
  XNOR2_X1 U478 ( .A(b[5]), .B(n320), .ZN(n222) );
  XNOR2_X1 U479 ( .A(b[4]), .B(n310), .ZN(n223) );
  XNOR2_X1 U480 ( .A(b[3]), .B(n313), .ZN(n224) );
  OAI22_X1 U481 ( .A1(n251), .A2(n259), .B1(n219), .B2(n342), .ZN(n167) );
  OAI22_X1 U482 ( .A1(n251), .A2(n218), .B1(n217), .B2(n342), .ZN(n184) );
  XNOR2_X1 U483 ( .A(b[6]), .B(n314), .ZN(n221) );
  INV_X1 U484 ( .A(n310), .ZN(n260) );
  XNOR2_X1 U485 ( .A(b[2]), .B(n320), .ZN(n225) );
  XNOR2_X1 U486 ( .A(b[7]), .B(n310), .ZN(n220) );
  XNOR2_X1 U487 ( .A(n313), .B(n351), .ZN(n227) );
  XNOR2_X1 U488 ( .A(b[1]), .B(n310), .ZN(n226) );
  XOR2_X1 U489 ( .A(n264), .B(a[2]), .Z(n248) );
  NAND2_X1 U490 ( .A1(n201), .A2(n169), .ZN(n97) );
  XNOR2_X1 U491 ( .A(b[5]), .B(n329), .ZN(n231) );
  XNOR2_X1 U492 ( .A(b[6]), .B(n329), .ZN(n230) );
  XNOR2_X1 U493 ( .A(b[4]), .B(n329), .ZN(n232) );
  XNOR2_X1 U494 ( .A(b[7]), .B(n316), .ZN(n229) );
  XNOR2_X1 U495 ( .A(b[3]), .B(n329), .ZN(n233) );
  XNOR2_X1 U496 ( .A(n329), .B(n351), .ZN(n236) );
  XNOR2_X1 U497 ( .A(b[2]), .B(n329), .ZN(n234) );
  XNOR2_X1 U498 ( .A(b[1]), .B(n329), .ZN(n235) );
  INV_X1 U499 ( .A(n316), .ZN(n261) );
  OAI21_X1 U500 ( .B1(n1), .B2(n19), .A(n20), .ZN(n18) );
  OAI21_X1 U501 ( .B1(n1), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X1 U502 ( .B1(n319), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U503 ( .B1(n319), .B2(n333), .A(n58), .ZN(n56) );
  OAI21_X1 U504 ( .B1(n319), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U505 ( .B1(n335), .B2(n64), .A(n65), .ZN(n63) );
  NAND2_X1 U506 ( .A1(n153), .A2(n168), .ZN(n89) );
  OAI22_X1 U507 ( .A1(n252), .A2(n221), .B1(n220), .B2(n347), .ZN(n128) );
  OAI22_X1 U508 ( .A1(n220), .A2(n252), .B1(n220), .B2(n347), .ZN(n160) );
  OAI22_X1 U509 ( .A1(n330), .A2(n222), .B1(n221), .B2(n347), .ZN(n187) );
  OAI22_X1 U510 ( .A1(n340), .A2(n224), .B1(n223), .B2(n347), .ZN(n189) );
  OAI22_X1 U511 ( .A1(n252), .A2(n225), .B1(n224), .B2(n347), .ZN(n190) );
  OAI22_X1 U512 ( .A1(n330), .A2(n223), .B1(n222), .B2(n347), .ZN(n188) );
  OAI22_X1 U513 ( .A1(n330), .A2(n260), .B1(n228), .B2(n347), .ZN(n168) );
  OAI22_X1 U514 ( .A1(n252), .A2(n226), .B1(n225), .B2(n347), .ZN(n191) );
  INV_X1 U515 ( .A(n347), .ZN(n161) );
  OAI22_X1 U516 ( .A1(n340), .A2(n227), .B1(n226), .B2(n347), .ZN(n192) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1_DW_mult_tc_2 ( a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50,
         n51, n52, n53, n56, n57, n58, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n80, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n92, n94, n95, n97, n98, n99, n100, n102,
         n103, n104, n105, n106, n108, n109, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n157, n160, n161, n163, n164, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n245, n246, n248, n249, n251, n252,
         n253, n254, n256, n258, n259, n260, n261, n262, n263, n264, n265,
         n273, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n351;
  assign n164 = a[0];
  assign n245 = b[0];
  assign n262 = a[7];
  assign n263 = a[5];
  assign n264 = a[3];
  assign n265 = a[1];

  FA_X1 U128 ( .A(n171), .B(n118), .CI(n178), .CO(n114), .S(n115) );
  FA_X1 U129 ( .A(n119), .B(n172), .CI(n122), .CO(n116), .S(n117) );
  FA_X1 U131 ( .A(n126), .B(n173), .CI(n123), .CO(n120), .S(n121) );
  FA_X1 U132 ( .A(n179), .B(n128), .CI(n186), .CO(n122), .S(n123) );
  FA_X1 U133 ( .A(n132), .B(n134), .CI(n127), .CO(n124), .S(n125) );
  FA_X1 U134 ( .A(n174), .B(n180), .CI(n129), .CO(n126), .S(n127) );
  FA_X1 U140 ( .A(n144), .B(n141), .CI(n139), .CO(n136), .S(n137) );
  FA_X1 U141 ( .A(n182), .B(n195), .CI(n188), .CO(n138), .S(n139) );
  HA_X1 U142 ( .A(n166), .B(n176), .CO(n140), .S(n141) );
  FA_X1 U144 ( .A(n196), .B(n177), .CI(n189), .CO(n144), .S(n145) );
  FA_X1 U145 ( .A(n190), .B(n197), .CI(n149), .CO(n146), .S(n147) );
  HA_X1 U146 ( .A(n167), .B(n184), .CO(n148), .S(n149) );
  FA_X1 U147 ( .A(n198), .B(n185), .CI(n191), .CO(n150), .S(n151) );
  HA_X1 U148 ( .A(n199), .B(n192), .CO(n152), .S(n153) );
  OR2_X2 U268 ( .A1(n339), .A2(n338), .ZN(n251) );
  XNOR2_X1 U269 ( .A(n303), .B(n133), .ZN(n131) );
  XNOR2_X1 U270 ( .A(n138), .B(n135), .ZN(n303) );
  OR2_X1 U271 ( .A1(n304), .A2(n338), .ZN(n326) );
  XOR2_X1 U272 ( .A(n264), .B(a[4]), .Z(n304) );
  INV_X1 U273 ( .A(n259), .ZN(n305) );
  CLKBUF_X1 U274 ( .A(n263), .Z(n306) );
  CLKBUF_X1 U275 ( .A(n340), .Z(n307) );
  BUF_X1 U276 ( .A(n265), .Z(n308) );
  INV_X1 U277 ( .A(n254), .ZN(n309) );
  XOR2_X1 U278 ( .A(n148), .B(n183), .Z(n310) );
  XOR2_X1 U279 ( .A(n145), .B(n310), .Z(n143) );
  NAND2_X1 U280 ( .A1(n145), .A2(n148), .ZN(n311) );
  NAND2_X1 U281 ( .A1(n145), .A2(n183), .ZN(n312) );
  NAND2_X1 U282 ( .A1(n148), .A2(n183), .ZN(n313) );
  NAND3_X1 U283 ( .A1(n311), .A2(n312), .A3(n313), .ZN(n142) );
  BUF_X1 U284 ( .A(n263), .Z(n330) );
  INV_X1 U285 ( .A(n341), .ZN(n314) );
  XNOR2_X1 U286 ( .A(n265), .B(n334), .ZN(n315) );
  NOR2_X1 U287 ( .A1(n64), .A2(n61), .ZN(n316) );
  NOR2_X2 U288 ( .A1(n121), .A2(n124), .ZN(n61) );
  OAI21_X1 U289 ( .B1(n61), .B2(n65), .A(n62), .ZN(n317) );
  NOR2_X2 U290 ( .A1(n131), .A2(n136), .ZN(n69) );
  XOR2_X1 U291 ( .A(n194), .B(n181), .Z(n318) );
  XOR2_X1 U292 ( .A(n318), .B(n140), .Z(n133) );
  NAND2_X1 U293 ( .A1(n194), .A2(n181), .ZN(n319) );
  NAND2_X1 U294 ( .A1(n194), .A2(n140), .ZN(n320) );
  NAND2_X1 U295 ( .A1(n181), .A2(n140), .ZN(n321) );
  NAND3_X1 U296 ( .A1(n319), .A2(n320), .A3(n321), .ZN(n132) );
  NAND2_X1 U297 ( .A1(n138), .A2(n135), .ZN(n322) );
  NAND2_X1 U298 ( .A1(n138), .A2(n133), .ZN(n323) );
  NAND2_X1 U299 ( .A1(n135), .A2(n133), .ZN(n324) );
  NAND3_X1 U300 ( .A1(n322), .A2(n323), .A3(n324), .ZN(n130) );
  INV_X1 U301 ( .A(n72), .ZN(n105) );
  OR2_X1 U302 ( .A1(n201), .A2(n169), .ZN(n325) );
  NAND2_X1 U303 ( .A1(n256), .A2(n248), .ZN(n327) );
  NAND2_X1 U304 ( .A1(n256), .A2(n248), .ZN(n252) );
  CLKBUF_X1 U305 ( .A(n264), .Z(n328) );
  CLKBUF_X1 U306 ( .A(n264), .Z(n329) );
  CLKBUF_X1 U307 ( .A(n264), .Z(n331) );
  XNOR2_X1 U308 ( .A(n330), .B(a[6]), .ZN(n332) );
  NAND2_X1 U309 ( .A1(n249), .A2(n273), .ZN(n333) );
  INV_X1 U310 ( .A(n164), .ZN(n334) );
  NAND2_X1 U311 ( .A1(n315), .A2(n273), .ZN(n253) );
  XOR2_X1 U312 ( .A(a[6]), .B(n262), .Z(n335) );
  OAI21_X2 U313 ( .B1(n84), .B2(n86), .A(n85), .ZN(n83) );
  BUF_X2 U314 ( .A(n245), .Z(n351) );
  XNOR2_X1 U315 ( .A(n265), .B(n334), .ZN(n249) );
  NAND2_X1 U316 ( .A1(n246), .A2(n254), .ZN(n336) );
  NAND2_X1 U317 ( .A1(n335), .A2(n254), .ZN(n337) );
  XNOR2_X1 U318 ( .A(n263), .B(a[4]), .ZN(n338) );
  XOR2_X1 U319 ( .A(n264), .B(a[4]), .Z(n339) );
  AOI21_X1 U320 ( .B1(n348), .B2(n83), .A(n80), .ZN(n340) );
  AOI21_X1 U321 ( .B1(n348), .B2(n83), .A(n80), .ZN(n78) );
  XNOR2_X2 U322 ( .A(n264), .B(a[4]), .ZN(n341) );
  OAI21_X1 U323 ( .B1(n76), .B2(n340), .A(n77), .ZN(n342) );
  XNOR2_X2 U324 ( .A(n265), .B(a[2]), .ZN(n343) );
  XNOR2_X1 U325 ( .A(n265), .B(a[2]), .ZN(n256) );
  AOI21_X1 U326 ( .B1(n67), .B2(n342), .A(n68), .ZN(n344) );
  AOI21_X1 U327 ( .B1(n67), .B2(n342), .A(n68), .ZN(n345) );
  AOI21_X1 U328 ( .B1(n67), .B2(n342), .A(n68), .ZN(n1) );
  XNOR2_X1 U329 ( .A(n263), .B(a[6]), .ZN(n346) );
  XNOR2_X1 U330 ( .A(n263), .B(a[6]), .ZN(n254) );
  XOR2_X1 U331 ( .A(n74), .B(n347), .Z(product[7]) );
  NAND2_X1 U332 ( .A1(n105), .A2(n73), .ZN(n347) );
  NOR2_X1 U333 ( .A1(n143), .A2(n146), .ZN(n76) );
  OR2_X1 U334 ( .A1(n147), .A2(n150), .ZN(n348) );
  NOR2_X1 U335 ( .A1(n151), .A2(n152), .ZN(n84) );
  INV_X2 U336 ( .A(n164), .ZN(n273) );
  INV_X1 U337 ( .A(n30), .ZN(n28) );
  INV_X1 U338 ( .A(n18), .ZN(product[15]) );
  OAI21_X1 U339 ( .B1(n344), .B2(n19), .A(n20), .ZN(n18) );
  NAND2_X1 U340 ( .A1(n103), .A2(n65), .ZN(n9) );
  INV_X1 U341 ( .A(n64), .ZN(n103) );
  INV_X1 U342 ( .A(n31), .ZN(n29) );
  NAND2_X1 U343 ( .A1(n52), .A2(n32), .ZN(n30) );
  NAND2_X1 U344 ( .A1(n348), .A2(n82), .ZN(n13) );
  NAND2_X1 U345 ( .A1(n102), .A2(n62), .ZN(n8) );
  XNOR2_X1 U346 ( .A(n16), .B(n95), .ZN(product[2]) );
  NAND2_X1 U347 ( .A1(n349), .A2(n94), .ZN(n16) );
  OAI21_X1 U348 ( .B1(n78), .B2(n76), .A(n77), .ZN(n75) );
  XNOR2_X1 U349 ( .A(n56), .B(n7), .ZN(product[11]) );
  NAND2_X1 U350 ( .A1(n52), .A2(n51), .ZN(n7) );
  XNOR2_X1 U351 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U352 ( .A1(n98), .A2(n24), .ZN(n4) );
  INV_X1 U353 ( .A(n23), .ZN(n98) );
  NAND2_X1 U354 ( .A1(n104), .A2(n70), .ZN(n10) );
  INV_X1 U355 ( .A(n82), .ZN(n80) );
  AOI21_X1 U356 ( .B1(n32), .B2(n53), .A(n33), .ZN(n31) );
  OAI21_X1 U357 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U358 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U359 ( .A1(n100), .A2(n44), .ZN(n6) );
  OAI21_X1 U360 ( .B1(n344), .B2(n46), .A(n47), .ZN(n45) );
  INV_X1 U361 ( .A(n50), .ZN(n52) );
  AOI21_X1 U362 ( .B1(n349), .B2(n95), .A(n92), .ZN(n90) );
  INV_X1 U363 ( .A(n94), .ZN(n92) );
  NOR2_X1 U364 ( .A1(n125), .A2(n130), .ZN(n64) );
  XNOR2_X1 U365 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U366 ( .A1(n99), .A2(n35), .ZN(n5) );
  OAI21_X1 U367 ( .B1(n344), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U368 ( .A(n34), .ZN(n99) );
  NAND2_X1 U369 ( .A1(n125), .A2(n130), .ZN(n65) );
  OAI21_X1 U370 ( .B1(n31), .B2(n23), .A(n24), .ZN(n22) );
  INV_X1 U371 ( .A(n51), .ZN(n53) );
  NOR2_X1 U372 ( .A1(n30), .A2(n23), .ZN(n21) );
  NAND2_X1 U373 ( .A1(n131), .A2(n136), .ZN(n70) );
  NAND2_X1 U374 ( .A1(n106), .A2(n77), .ZN(n12) );
  INV_X1 U375 ( .A(n76), .ZN(n106) );
  XOR2_X1 U376 ( .A(n15), .B(n90), .Z(product[3]) );
  INV_X1 U377 ( .A(n88), .ZN(n109) );
  OR2_X1 U378 ( .A1(n187), .A2(n175), .ZN(n134) );
  NOR2_X1 U379 ( .A1(n170), .A2(n112), .ZN(n23) );
  NOR2_X1 U380 ( .A1(n116), .A2(n115), .ZN(n41) );
  INV_X1 U381 ( .A(n112), .ZN(n113) );
  XNOR2_X1 U382 ( .A(n187), .B(n175), .ZN(n135) );
  NAND2_X1 U383 ( .A1(n116), .A2(n115), .ZN(n44) );
  NOR2_X1 U384 ( .A1(n114), .A2(n113), .ZN(n34) );
  NAND2_X1 U385 ( .A1(n170), .A2(n112), .ZN(n24) );
  INV_X1 U386 ( .A(n97), .ZN(n95) );
  NOR2_X1 U387 ( .A1(n137), .A2(n142), .ZN(n72) );
  OR2_X1 U388 ( .A1(n200), .A2(n193), .ZN(n349) );
  NOR2_X1 U389 ( .A1(n117), .A2(n120), .ZN(n50) );
  INV_X1 U390 ( .A(n87), .ZN(n86) );
  NAND2_X1 U391 ( .A1(n114), .A2(n113), .ZN(n35) );
  NAND2_X1 U392 ( .A1(n117), .A2(n120), .ZN(n51) );
  NAND2_X1 U393 ( .A1(n137), .A2(n142), .ZN(n73) );
  NAND2_X1 U394 ( .A1(n143), .A2(n146), .ZN(n77) );
  NAND2_X1 U395 ( .A1(n121), .A2(n124), .ZN(n62) );
  XOR2_X1 U396 ( .A(n14), .B(n86), .Z(product[4]) );
  NAND2_X1 U397 ( .A1(n108), .A2(n85), .ZN(n14) );
  INV_X1 U398 ( .A(n84), .ZN(n108) );
  AND2_X1 U399 ( .A1(n351), .A2(n309), .ZN(n177) );
  INV_X1 U400 ( .A(n118), .ZN(n119) );
  AND2_X1 U401 ( .A1(n351), .A2(n314), .ZN(n185) );
  INV_X1 U402 ( .A(n157), .ZN(n178) );
  OR2_X1 U403 ( .A1(n351), .A2(n259), .ZN(n219) );
  AND2_X1 U404 ( .A1(n325), .A2(n97), .ZN(product[1]) );
  INV_X1 U405 ( .A(n163), .ZN(n194) );
  INV_X1 U406 ( .A(n128), .ZN(n129) );
  NAND2_X1 U407 ( .A1(n151), .A2(n152), .ZN(n85) );
  INV_X1 U408 ( .A(n154), .ZN(n170) );
  OR2_X1 U409 ( .A1(n351), .A2(n258), .ZN(n210) );
  INV_X1 U410 ( .A(n160), .ZN(n186) );
  AND2_X1 U411 ( .A1(n351), .A2(n161), .ZN(n193) );
  OR2_X1 U412 ( .A1(n351), .A2(n260), .ZN(n228) );
  OR2_X1 U413 ( .A1(n351), .A2(n261), .ZN(n237) );
  XNOR2_X1 U414 ( .A(b[4]), .B(n262), .ZN(n205) );
  XNOR2_X1 U415 ( .A(b[7]), .B(n262), .ZN(n202) );
  XNOR2_X1 U416 ( .A(b[5]), .B(n262), .ZN(n204) );
  XNOR2_X1 U417 ( .A(b[6]), .B(n262), .ZN(n203) );
  XOR2_X1 U418 ( .A(a[6]), .B(n262), .Z(n246) );
  XNOR2_X1 U419 ( .A(n262), .B(n351), .ZN(n209) );
  INV_X1 U420 ( .A(n262), .ZN(n258) );
  AND2_X1 U421 ( .A1(n351), .A2(n164), .ZN(product[0]) );
  OAI21_X1 U422 ( .B1(n26), .B2(n345), .A(n27), .ZN(n25) );
  OAI21_X1 U423 ( .B1(n345), .B2(n57), .A(n58), .ZN(n56) );
  NAND2_X1 U424 ( .A1(n147), .A2(n150), .ZN(n82) );
  AOI21_X1 U425 ( .B1(n317), .B2(n21), .A(n22), .ZN(n20) );
  AOI21_X1 U426 ( .B1(n317), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U427 ( .B1(n2), .B2(n52), .A(n53), .ZN(n47) );
  INV_X1 U428 ( .A(n317), .ZN(n58) );
  INV_X1 U429 ( .A(n61), .ZN(n102) );
  AOI21_X1 U430 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  NOR2_X1 U431 ( .A1(n64), .A2(n61), .ZN(n3) );
  OAI21_X1 U432 ( .B1(n61), .B2(n65), .A(n62), .ZN(n2) );
  XNOR2_X1 U433 ( .A(n71), .B(n10), .ZN(product[8]) );
  XNOR2_X1 U434 ( .A(n13), .B(n83), .ZN(product[5]) );
  OAI22_X1 U435 ( .A1(n333), .A2(n232), .B1(n231), .B2(n273), .ZN(n197) );
  OAI22_X1 U436 ( .A1(n333), .A2(n231), .B1(n230), .B2(n273), .ZN(n196) );
  OAI22_X1 U437 ( .A1(n253), .A2(n234), .B1(n233), .B2(n273), .ZN(n199) );
  OAI22_X1 U438 ( .A1(n333), .A2(n233), .B1(n232), .B2(n273), .ZN(n198) );
  OAI22_X1 U439 ( .A1(n333), .A2(n235), .B1(n234), .B2(n273), .ZN(n200) );
  OAI22_X1 U440 ( .A1(n253), .A2(n261), .B1(n237), .B2(n273), .ZN(n169) );
  NAND2_X1 U441 ( .A1(n316), .A2(n21), .ZN(n19) );
  NAND2_X1 U442 ( .A1(n316), .A2(n28), .ZN(n26) );
  NAND2_X1 U443 ( .A1(n316), .A2(n39), .ZN(n37) );
  INV_X1 U444 ( .A(n3), .ZN(n57) );
  NAND2_X1 U445 ( .A1(n3), .A2(n52), .ZN(n46) );
  NOR2_X1 U446 ( .A1(n41), .A2(n34), .ZN(n32) );
  INV_X1 U447 ( .A(n41), .ZN(n100) );
  NOR2_X1 U448 ( .A1(n50), .A2(n41), .ZN(n39) );
  OAI21_X1 U449 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  INV_X1 U450 ( .A(n69), .ZN(n104) );
  NOR2_X1 U451 ( .A1(n69), .A2(n72), .ZN(n67) );
  OAI21_X1 U452 ( .B1(n69), .B2(n73), .A(n70), .ZN(n68) );
  XOR2_X1 U453 ( .A(n345), .B(n9), .Z(product[9]) );
  OAI22_X1 U454 ( .A1(n253), .A2(n236), .B1(n235), .B2(n273), .ZN(n201) );
  OAI21_X1 U455 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  INV_X1 U456 ( .A(n329), .ZN(n260) );
  XNOR2_X1 U457 ( .A(n331), .B(b[5]), .ZN(n222) );
  XNOR2_X1 U458 ( .A(n328), .B(n351), .ZN(n227) );
  XNOR2_X1 U459 ( .A(n328), .B(b[4]), .ZN(n223) );
  XNOR2_X1 U460 ( .A(n331), .B(b[6]), .ZN(n221) );
  XOR2_X1 U461 ( .A(n264), .B(a[2]), .Z(n248) );
  OAI22_X1 U462 ( .A1(n333), .A2(n230), .B1(n229), .B2(n273), .ZN(n195) );
  OAI22_X1 U463 ( .A1(n229), .A2(n253), .B1(n229), .B2(n273), .ZN(n163) );
  XOR2_X1 U464 ( .A(n12), .B(n307), .Z(product[6]) );
  XNOR2_X1 U465 ( .A(n329), .B(b[7]), .ZN(n220) );
  NAND2_X1 U466 ( .A1(n109), .A2(n89), .ZN(n15) );
  OAI21_X1 U467 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  XNOR2_X1 U468 ( .A(b[3]), .B(n262), .ZN(n206) );
  XNOR2_X1 U469 ( .A(n329), .B(b[3]), .ZN(n224) );
  NAND2_X1 U470 ( .A1(n200), .A2(n193), .ZN(n94) );
  XNOR2_X1 U471 ( .A(b[2]), .B(n262), .ZN(n207) );
  XNOR2_X1 U472 ( .A(n331), .B(b[2]), .ZN(n225) );
  XNOR2_X1 U473 ( .A(n328), .B(b[1]), .ZN(n226) );
  XNOR2_X1 U474 ( .A(b[1]), .B(n262), .ZN(n208) );
  NAND2_X1 U475 ( .A1(n153), .A2(n168), .ZN(n89) );
  NOR2_X1 U476 ( .A1(n153), .A2(n168), .ZN(n88) );
  XNOR2_X1 U477 ( .A(n308), .B(b[5]), .ZN(n231) );
  XNOR2_X1 U478 ( .A(n265), .B(b[6]), .ZN(n230) );
  XNOR2_X1 U479 ( .A(n308), .B(b[4]), .ZN(n232) );
  XNOR2_X1 U480 ( .A(n308), .B(n351), .ZN(n236) );
  INV_X1 U481 ( .A(n265), .ZN(n261) );
  XNOR2_X1 U482 ( .A(n265), .B(b[7]), .ZN(n229) );
  XNOR2_X1 U483 ( .A(n265), .B(b[1]), .ZN(n235) );
  XNOR2_X1 U484 ( .A(n265), .B(b[2]), .ZN(n234) );
  XNOR2_X1 U485 ( .A(n265), .B(b[3]), .ZN(n233) );
  OAI22_X1 U486 ( .A1(n326), .A2(n217), .B1(n216), .B2(n341), .ZN(n183) );
  OAI22_X1 U487 ( .A1(n326), .A2(n212), .B1(n211), .B2(n341), .ZN(n118) );
  OAI22_X1 U488 ( .A1(n211), .A2(n326), .B1(n211), .B2(n341), .ZN(n157) );
  OAI22_X1 U489 ( .A1(n326), .A2(n213), .B1(n212), .B2(n341), .ZN(n179) );
  OAI22_X1 U490 ( .A1(n326), .A2(n214), .B1(n213), .B2(n341), .ZN(n180) );
  OAI22_X1 U491 ( .A1(n326), .A2(n216), .B1(n215), .B2(n341), .ZN(n182) );
  OAI22_X1 U492 ( .A1(n251), .A2(n215), .B1(n214), .B2(n341), .ZN(n181) );
  OAI22_X1 U493 ( .A1(n251), .A2(n259), .B1(n219), .B2(n341), .ZN(n167) );
  OAI22_X1 U494 ( .A1(n251), .A2(n218), .B1(n217), .B2(n341), .ZN(n184) );
  INV_X1 U495 ( .A(n75), .ZN(n74) );
  NAND2_X1 U496 ( .A1(n201), .A2(n169), .ZN(n97) );
  OAI22_X1 U497 ( .A1(n202), .A2(n336), .B1(n202), .B2(n332), .ZN(n154) );
  OAI22_X1 U498 ( .A1(n336), .A2(n206), .B1(n346), .B2(n205), .ZN(n173) );
  OAI22_X1 U499 ( .A1(n337), .A2(n203), .B1(n332), .B2(n202), .ZN(n112) );
  OAI22_X1 U500 ( .A1(n336), .A2(n205), .B1(n332), .B2(n204), .ZN(n172) );
  OAI22_X1 U501 ( .A1(n337), .A2(n204), .B1(n346), .B2(n203), .ZN(n171) );
  OAI22_X1 U502 ( .A1(n337), .A2(n208), .B1(n346), .B2(n207), .ZN(n175) );
  OAI22_X1 U503 ( .A1(n336), .A2(n207), .B1(n346), .B2(n206), .ZN(n174) );
  XNOR2_X1 U504 ( .A(n330), .B(b[7]), .ZN(n211) );
  OAI22_X1 U505 ( .A1(n336), .A2(n258), .B1(n210), .B2(n346), .ZN(n166) );
  OAI22_X1 U506 ( .A1(n337), .A2(n209), .B1(n346), .B2(n208), .ZN(n176) );
  XNOR2_X1 U507 ( .A(n330), .B(b[6]), .ZN(n212) );
  XNOR2_X1 U508 ( .A(n306), .B(b[5]), .ZN(n213) );
  XNOR2_X1 U509 ( .A(n306), .B(b[2]), .ZN(n216) );
  XNOR2_X1 U510 ( .A(n305), .B(b[3]), .ZN(n215) );
  XNOR2_X1 U511 ( .A(n263), .B(b[4]), .ZN(n214) );
  XNOR2_X1 U512 ( .A(n305), .B(n351), .ZN(n218) );
  INV_X1 U513 ( .A(n263), .ZN(n259) );
  XNOR2_X1 U514 ( .A(n263), .B(b[1]), .ZN(n217) );
  XNOR2_X1 U515 ( .A(n63), .B(n8), .ZN(product[10]) );
  OAI21_X1 U516 ( .B1(n1), .B2(n64), .A(n65), .ZN(n63) );
  OAI22_X1 U517 ( .A1(n327), .A2(n221), .B1(n220), .B2(n343), .ZN(n128) );
  OAI22_X1 U518 ( .A1(n220), .A2(n252), .B1(n220), .B2(n343), .ZN(n160) );
  OAI22_X1 U519 ( .A1(n327), .A2(n222), .B1(n221), .B2(n343), .ZN(n187) );
  OAI22_X1 U520 ( .A1(n252), .A2(n224), .B1(n223), .B2(n343), .ZN(n189) );
  OAI22_X1 U521 ( .A1(n327), .A2(n225), .B1(n224), .B2(n343), .ZN(n190) );
  OAI22_X1 U522 ( .A1(n327), .A2(n223), .B1(n222), .B2(n343), .ZN(n188) );
  OAI22_X1 U523 ( .A1(n327), .A2(n260), .B1(n228), .B2(n343), .ZN(n168) );
  OAI22_X1 U524 ( .A1(n327), .A2(n226), .B1(n225), .B2(n343), .ZN(n191) );
  INV_X1 U525 ( .A(n343), .ZN(n161) );
  OAI22_X1 U526 ( .A1(n252), .A2(n227), .B1(n226), .B2(n343), .ZN(n192) );
endmodule


module mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1 ( ia, ix, out );
  input [7:0] ia;
  input [7:0] ix;
  output [15:0] out;


  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1_DW_mult_tc_2 mult_44 ( .a(ia), .b(
        ix), .product(out) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_1_DW01_add_2 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n8, n10, n11, n12, n13, n14, n15, n16, n19, n20,
         n21, n22, n24, n26, n27, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n51, n52, n54, n56,
         n57, n58, n60, n62, n63, n64, n65, n66, n68, n70, n71, n72, n73, n74,
         n76, n78, n79, n80, n81, n82, n84, n86, n87, n89, n92, n93, n95, n99,
         n101, n103, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188;

  OR2_X2 U125 ( .A1(A[14]), .A2(B[14]), .ZN(n184) );
  AOI21_X1 U126 ( .B1(n71), .B2(n168), .A(n68), .ZN(n160) );
  BUF_X1 U127 ( .A(n40), .Z(n161) );
  NOR2_X1 U128 ( .A1(B[12]), .A2(A[12]), .ZN(n35) );
  CLKBUF_X1 U129 ( .A(n178), .Z(n162) );
  CLKBUF_X1 U130 ( .A(n43), .Z(n163) );
  CLKBUF_X1 U131 ( .A(B[11]), .Z(n164) );
  BUF_X1 U132 ( .A(n36), .Z(n165) );
  BUF_X1 U133 ( .A(n33), .Z(n166) );
  CLKBUF_X1 U134 ( .A(A[11]), .Z(n167) );
  OR2_X1 U135 ( .A1(B[5]), .A2(A[5]), .ZN(n168) );
  OR2_X1 U136 ( .A1(B[15]), .A2(A[15]), .ZN(n169) );
  OR2_X1 U137 ( .A1(B[0]), .A2(A[0]), .ZN(n170) );
  AND2_X1 U138 ( .A1(n170), .A2(n89), .ZN(SUM[0]) );
  XNOR2_X1 U139 ( .A(n44), .B(n172), .ZN(SUM[10]) );
  AND2_X1 U140 ( .A1(n95), .A2(n43), .ZN(n172) );
  XNOR2_X1 U141 ( .A(n41), .B(n173), .ZN(SUM[11]) );
  NAND2_X1 U142 ( .A1(n177), .A2(n161), .ZN(n173) );
  OR2_X1 U143 ( .A1(A[9]), .A2(B[9]), .ZN(n174) );
  OR2_X1 U144 ( .A1(B[9]), .A2(A[9]), .ZN(n182) );
  INV_X1 U145 ( .A(n95), .ZN(n175) );
  NOR2_X1 U146 ( .A1(A[11]), .A2(B[11]), .ZN(n176) );
  INV_X1 U147 ( .A(n180), .ZN(n51) );
  OR2_X1 U148 ( .A1(n164), .A2(n167), .ZN(n177) );
  NOR2_X1 U149 ( .A1(A[11]), .A2(B[11]), .ZN(n39) );
  NOR2_X1 U150 ( .A1(B[13]), .A2(A[13]), .ZN(n178) );
  OR2_X1 U151 ( .A1(n178), .A2(n35), .ZN(n179) );
  AND2_X1 U152 ( .A1(B[9]), .A2(A[9]), .ZN(n180) );
  XNOR2_X1 U153 ( .A(n181), .B(n57), .ZN(SUM[8]) );
  NAND2_X1 U154 ( .A1(n183), .A2(n56), .ZN(n181) );
  INV_X1 U155 ( .A(n58), .ZN(n57) );
  INV_X1 U156 ( .A(n62), .ZN(n60) );
  AOI21_X1 U157 ( .B1(n71), .B2(n168), .A(n68), .ZN(n66) );
  INV_X1 U158 ( .A(n70), .ZN(n68) );
  INV_X1 U159 ( .A(n42), .ZN(n95) );
  NAND2_X1 U160 ( .A1(n93), .A2(n165), .ZN(n5) );
  OAI21_X1 U161 ( .B1(n64), .B2(n66), .A(n65), .ZN(n63) );
  XOR2_X1 U162 ( .A(n8), .B(n52), .Z(SUM[9]) );
  AOI21_X1 U163 ( .B1(n183), .B2(n57), .A(n54), .ZN(n52) );
  XNOR2_X1 U164 ( .A(n12), .B(n71), .ZN(SUM[5]) );
  NAND2_X1 U165 ( .A1(n168), .A2(n70), .ZN(n12) );
  NAND2_X1 U166 ( .A1(n99), .A2(n65), .ZN(n11) );
  INV_X1 U167 ( .A(n64), .ZN(n99) );
  NAND2_X1 U168 ( .A1(n92), .A2(n166), .ZN(n4) );
  NAND2_X1 U169 ( .A1(n185), .A2(n62), .ZN(n10) );
  OAI21_X1 U170 ( .B1(n72), .B2(n74), .A(n73), .ZN(n71) );
  OR2_X1 U171 ( .A1(B[8]), .A2(A[8]), .ZN(n183) );
  NOR2_X1 U172 ( .A1(A[10]), .A2(B[10]), .ZN(n42) );
  AOI21_X1 U173 ( .B1(n186), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U174 ( .A(n78), .ZN(n76) );
  NAND2_X1 U175 ( .A1(B[12]), .A2(A[12]), .ZN(n36) );
  XOR2_X1 U176 ( .A(n13), .B(n74), .Z(SUM[4]) );
  NAND2_X1 U177 ( .A1(n101), .A2(n73), .ZN(n13) );
  INV_X1 U178 ( .A(n72), .ZN(n101) );
  NOR2_X1 U179 ( .A1(B[6]), .A2(A[6]), .ZN(n64) );
  NAND2_X1 U180 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  NAND2_X1 U181 ( .A1(B[6]), .A2(A[6]), .ZN(n65) );
  XNOR2_X1 U182 ( .A(n14), .B(n79), .ZN(SUM[3]) );
  NAND2_X1 U183 ( .A1(n186), .A2(n78), .ZN(n14) );
  OR2_X1 U184 ( .A1(B[7]), .A2(A[7]), .ZN(n185) );
  NAND2_X1 U185 ( .A1(n169), .A2(n19), .ZN(n2) );
  OAI21_X1 U186 ( .B1(n82), .B2(n80), .A(n81), .ZN(n79) );
  OR2_X1 U187 ( .A1(B[3]), .A2(A[3]), .ZN(n186) );
  NOR2_X1 U188 ( .A1(B[4]), .A2(A[4]), .ZN(n72) );
  NAND2_X1 U189 ( .A1(B[4]), .A2(A[4]), .ZN(n73) );
  NAND2_X1 U190 ( .A1(n103), .A2(n81), .ZN(n15) );
  INV_X1 U191 ( .A(n80), .ZN(n103) );
  AOI21_X1 U192 ( .B1(n187), .B2(n87), .A(n84), .ZN(n82) );
  INV_X1 U193 ( .A(n86), .ZN(n84) );
  NOR2_X1 U194 ( .A1(B[2]), .A2(A[2]), .ZN(n80) );
  NAND2_X1 U195 ( .A1(B[2]), .A2(A[2]), .ZN(n81) );
  NAND2_X1 U196 ( .A1(n187), .A2(n86), .ZN(n16) );
  INV_X1 U197 ( .A(n89), .ZN(n87) );
  NAND2_X1 U198 ( .A1(B[1]), .A2(A[1]), .ZN(n86) );
  OR2_X1 U199 ( .A1(B[1]), .A2(A[1]), .ZN(n187) );
  NAND2_X1 U200 ( .A1(B[0]), .A2(A[0]), .ZN(n89) );
  XOR2_X1 U201 ( .A(n15), .B(n82), .Z(SUM[2]) );
  XNOR2_X1 U202 ( .A(n16), .B(n87), .ZN(SUM[1]) );
  AOI21_X1 U203 ( .B1(n45), .B2(n37), .A(n38), .ZN(n188) );
  AOI21_X1 U204 ( .B1(n45), .B2(n37), .A(n38), .ZN(n1) );
  NOR2_X1 U205 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  XNOR2_X1 U206 ( .A(n10), .B(n63), .ZN(SUM[7]) );
  AOI21_X1 U207 ( .B1(n63), .B2(n185), .A(n60), .ZN(n58) );
  NAND2_X1 U208 ( .A1(B[5]), .A2(A[5]), .ZN(n70) );
  INV_X1 U209 ( .A(n26), .ZN(n24) );
  NAND2_X1 U210 ( .A1(n184), .A2(n26), .ZN(n3) );
  AOI21_X1 U211 ( .B1(n182), .B2(n54), .A(n180), .ZN(n47) );
  XOR2_X1 U212 ( .A(n11), .B(n160), .Z(SUM[6]) );
  NAND2_X1 U213 ( .A1(B[3]), .A2(A[3]), .ZN(n78) );
  INV_X1 U214 ( .A(n56), .ZN(n54) );
  NAND2_X1 U215 ( .A1(B[8]), .A2(A[8]), .ZN(n56) );
  NAND2_X1 U216 ( .A1(B[11]), .A2(A[11]), .ZN(n40) );
  NAND2_X1 U217 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NAND2_X1 U218 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  INV_X1 U219 ( .A(n162), .ZN(n92) );
  NOR2_X1 U220 ( .A1(n178), .A2(n35), .ZN(n30) );
  OAI21_X1 U221 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  NAND2_X1 U222 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  NAND2_X1 U223 ( .A1(A[10]), .A2(B[10]), .ZN(n43) );
  NAND2_X1 U224 ( .A1(n30), .A2(n184), .ZN(n21) );
  OAI21_X1 U225 ( .B1(n39), .B2(n43), .A(n40), .ZN(n38) );
  NOR2_X1 U226 ( .A1(n176), .A2(n42), .ZN(n37) );
  OAI21_X1 U227 ( .B1(n44), .B2(n175), .A(n163), .ZN(n41) );
  XNOR2_X1 U228 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  INV_X1 U229 ( .A(n45), .ZN(n44) );
  INV_X1 U230 ( .A(n35), .ZN(n93) );
  AOI21_X1 U231 ( .B1(n31), .B2(n184), .A(n24), .ZN(n22) );
  INV_X1 U232 ( .A(n31), .ZN(n29) );
  XNOR2_X1 U233 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  OAI21_X1 U234 ( .B1(n46), .B2(n58), .A(n47), .ZN(n45) );
  XNOR2_X1 U235 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XOR2_X1 U236 ( .A(n188), .B(n5), .Z(SUM[12]) );
  OAI21_X1 U237 ( .B1(n21), .B2(n1), .A(n22), .ZN(n20) );
  OAI21_X1 U238 ( .B1(n188), .B2(n179), .A(n29), .ZN(n27) );
  OAI21_X1 U239 ( .B1(n1), .B2(n35), .A(n165), .ZN(n34) );
  NAND2_X1 U240 ( .A1(n51), .A2(n174), .ZN(n8) );
  NAND2_X1 U241 ( .A1(n174), .A2(n183), .ZN(n46) );
endmodule


module recursive_add_layer_INPUT_SCALE2_WIDTH16_1 ( .in({\in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] ,
         \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] ,
         \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] ,
         \in[1][0] , \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] ,
         \in[0][11] , \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] ,
         \in[0][6] , \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] ,
         \in[0][1] , \in[0][0] ;


  recursive_add_layer_INPUT_SCALE2_WIDTH16_1_DW01_add_2 add_56 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM(out) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_1_DW01_add_4 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n9, n12, n13, n14, n15, n16, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n59, n60, n62, n64, n65, n66, n68, n70, n71, n72, n73,
         n74, n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89, n91, n93,
         n94, n95, n97, n98, n102, n104, n106, n162, n163, n164, n165, n166,
         n167, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183;

  OR2_X1 U127 ( .A1(B[11]), .A2(A[11]), .ZN(n162) );
  CLKBUF_X1 U128 ( .A(n51), .Z(n163) );
  OR2_X1 U129 ( .A1(B[8]), .A2(A[8]), .ZN(n164) );
  OR2_X1 U130 ( .A1(B[8]), .A2(A[8]), .ZN(n181) );
  INV_X1 U131 ( .A(n165), .ZN(n59) );
  AND2_X1 U132 ( .A1(B[8]), .A2(A[8]), .ZN(n165) );
  INV_X1 U133 ( .A(n36), .ZN(n166) );
  NOR2_X1 U134 ( .A1(A[12]), .A2(B[12]), .ZN(n167) );
  NOR2_X1 U135 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  AND2_X1 U136 ( .A1(n170), .A2(n91), .ZN(SUM[0]) );
  OR2_X1 U137 ( .A1(B[6]), .A2(A[6]), .ZN(n169) );
  OR2_X1 U138 ( .A1(B[0]), .A2(A[0]), .ZN(n170) );
  INV_X1 U139 ( .A(n98), .ZN(n171) );
  CLKBUF_X1 U140 ( .A(n1), .Z(n172) );
  XNOR2_X1 U141 ( .A(n1), .B(n173), .ZN(SUM[11]) );
  AND2_X1 U142 ( .A1(n162), .A2(n43), .ZN(n173) );
  NOR2_X1 U143 ( .A1(A[10]), .A2(B[10]), .ZN(n174) );
  NOR2_X1 U144 ( .A1(A[10]), .A2(B[10]), .ZN(n47) );
  INV_X1 U145 ( .A(n50), .ZN(n98) );
  XOR2_X1 U146 ( .A(n175), .B(n71), .Z(SUM[6]) );
  AND2_X1 U147 ( .A1(n169), .A2(n70), .ZN(n175) );
  XOR2_X1 U148 ( .A(n176), .B(n65), .Z(SUM[7]) );
  AND2_X1 U149 ( .A1(n180), .A2(n64), .ZN(n176) );
  XOR2_X1 U150 ( .A(n49), .B(n177), .Z(SUM[10]) );
  AND2_X1 U151 ( .A1(n97), .A2(n48), .ZN(n177) );
  AOI21_X2 U152 ( .B1(n53), .B2(n45), .A(n46), .ZN(n1) );
  OR2_X1 U153 ( .A1(B[7]), .A2(A[7]), .ZN(n180) );
  XNOR2_X1 U154 ( .A(n52), .B(n178), .ZN(SUM[9]) );
  AND2_X1 U155 ( .A1(n98), .A2(n51), .ZN(n178) );
  INV_X1 U156 ( .A(n66), .ZN(n65) );
  OAI21_X1 U157 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  AOI21_X1 U158 ( .B1(n169), .B2(n71), .A(n68), .ZN(n66) );
  INV_X1 U159 ( .A(n70), .ZN(n68) );
  OAI21_X1 U160 ( .B1(n167), .B2(n43), .A(n40), .ZN(n38) );
  OAI21_X1 U161 ( .B1(n54), .B2(n66), .A(n55), .ZN(n53) );
  AOI21_X1 U162 ( .B1(n181), .B2(n62), .A(n165), .ZN(n55) );
  XOR2_X1 U163 ( .A(n60), .B(n9), .Z(SUM[8]) );
  AOI21_X1 U164 ( .B1(n65), .B2(n180), .A(n62), .ZN(n60) );
  INV_X1 U165 ( .A(n33), .ZN(n31) );
  NAND2_X1 U166 ( .A1(n95), .A2(n40), .ZN(n5) );
  NAND2_X1 U167 ( .A1(n179), .A2(n19), .ZN(n2) );
  NAND2_X1 U168 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NOR2_X1 U169 ( .A1(n42), .A2(n39), .ZN(n37) );
  XNOR2_X1 U170 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U171 ( .A1(n93), .A2(n26), .ZN(n3) );
  INV_X1 U172 ( .A(n25), .ZN(n93) );
  INV_X1 U173 ( .A(n64), .ZN(n62) );
  OAI21_X1 U174 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  NOR2_X1 U175 ( .A1(n32), .A2(n25), .ZN(n23) );
  OR2_X1 U176 ( .A1(B[15]), .A2(A[15]), .ZN(n179) );
  INV_X1 U177 ( .A(n32), .ZN(n94) );
  NAND2_X1 U178 ( .A1(n102), .A2(n73), .ZN(n12) );
  INV_X1 U179 ( .A(n72), .ZN(n102) );
  NOR2_X1 U180 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  INV_X1 U181 ( .A(n78), .ZN(n76) );
  XOR2_X1 U182 ( .A(n14), .B(n82), .Z(SUM[3]) );
  NAND2_X1 U183 ( .A1(n104), .A2(n81), .ZN(n14) );
  INV_X1 U184 ( .A(n80), .ZN(n104) );
  NOR2_X1 U185 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND2_X1 U186 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  OAI21_X1 U187 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  NOR2_X1 U188 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  OR2_X1 U189 ( .A1(B[2]), .A2(A[2]), .ZN(n182) );
  NAND2_X1 U190 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
  NAND2_X1 U191 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  NAND2_X1 U192 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  NAND2_X1 U193 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U194 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  XNOR2_X1 U195 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  NAND2_X1 U196 ( .A1(n183), .A2(n78), .ZN(n13) );
  XNOR2_X1 U197 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U198 ( .A1(n182), .A2(n86), .ZN(n15) );
  AOI21_X1 U199 ( .B1(n87), .B2(n182), .A(n84), .ZN(n82) );
  INV_X1 U200 ( .A(n86), .ZN(n84) );
  NOR2_X1 U201 ( .A1(B[3]), .A2(A[3]), .ZN(n80) );
  OR2_X1 U202 ( .A1(B[4]), .A2(A[4]), .ZN(n183) );
  NAND2_X1 U203 ( .A1(B[3]), .A2(A[3]), .ZN(n81) );
  NAND2_X1 U204 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  XOR2_X1 U205 ( .A(n16), .B(n91), .Z(SUM[1]) );
  NAND2_X1 U206 ( .A1(n106), .A2(n89), .ZN(n16) );
  INV_X1 U207 ( .A(n88), .ZN(n106) );
  OAI21_X1 U208 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U209 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U210 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  NAND2_X1 U211 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  NAND2_X1 U212 ( .A1(n94), .A2(n33), .ZN(n4) );
  NAND2_X1 U213 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  NAND2_X1 U214 ( .A1(A[12]), .A2(B[12]), .ZN(n40) );
  XNOR2_X1 U215 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  NAND2_X1 U216 ( .A1(A[9]), .A2(B[9]), .ZN(n51) );
  XNOR2_X1 U217 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  XNOR2_X1 U218 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  XOR2_X1 U219 ( .A(n12), .B(n74), .Z(SUM[5]) );
  AOI21_X1 U220 ( .B1(n183), .B2(n79), .A(n76), .ZN(n74) );
  NOR2_X1 U221 ( .A1(B[11]), .A2(A[11]), .ZN(n42) );
  NAND2_X1 U222 ( .A1(n37), .A2(n23), .ZN(n21) );
  INV_X1 U223 ( .A(n37), .ZN(n35) );
  NAND2_X1 U224 ( .A1(n37), .A2(n94), .ZN(n28) );
  NOR2_X1 U225 ( .A1(B[9]), .A2(A[9]), .ZN(n50) );
  INV_X1 U226 ( .A(n174), .ZN(n97) );
  NOR2_X1 U227 ( .A1(n174), .A2(n50), .ZN(n45) );
  OAI21_X1 U228 ( .B1(n47), .B2(n51), .A(n48), .ZN(n46) );
  INV_X1 U229 ( .A(n38), .ZN(n36) );
  AOI21_X1 U230 ( .B1(n166), .B2(n23), .A(n24), .ZN(n22) );
  AOI21_X1 U231 ( .B1(n38), .B2(n94), .A(n31), .ZN(n29) );
  INV_X1 U232 ( .A(n167), .ZN(n95) );
  OAI21_X1 U233 ( .B1(n52), .B2(n171), .A(n163), .ZN(n49) );
  NAND2_X1 U234 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  INV_X1 U235 ( .A(n53), .ZN(n52) );
  OAI21_X1 U236 ( .B1(n172), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U237 ( .B1(n28), .B2(n1), .A(n29), .ZN(n27) );
  OAI21_X1 U238 ( .B1(n1), .B2(n35), .A(n36), .ZN(n34) );
  OAI21_X1 U239 ( .B1(n1), .B2(n42), .A(n43), .ZN(n41) );
  NAND2_X1 U240 ( .A1(n164), .A2(n59), .ZN(n9) );
  NAND2_X1 U241 ( .A1(n164), .A2(n180), .ZN(n54) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_1_DW01_add_5 ( A, B, CI, SUM, 
        CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n9, n10, n12, n13, n14, n15, n16, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n59, n60, n62, n64, n65, n66, n68, n70, n71, n72, n73, n74,
         n76, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89, n91, n93, n95,
         n97, n98, n102, n104, n106, n162, n163, n164, n165, n166, n167, n168,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187;

  AOI21_X1 U127 ( .B1(n186), .B2(n62), .A(n174), .ZN(n162) );
  BUF_X1 U128 ( .A(n47), .Z(n163) );
  OAI21_X1 U129 ( .B1(n54), .B2(n66), .A(n162), .ZN(n164) );
  OAI21_X1 U130 ( .B1(n54), .B2(n66), .A(n55), .ZN(n53) );
  OR2_X1 U131 ( .A1(n42), .A2(n168), .ZN(n165) );
  OR2_X1 U132 ( .A1(B[13]), .A2(A[13]), .ZN(n166) );
  CLKBUF_X1 U133 ( .A(n1), .Z(n167) );
  NOR2_X1 U134 ( .A1(B[12]), .A2(A[12]), .ZN(n168) );
  NOR2_X1 U135 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  INV_X1 U136 ( .A(n174), .ZN(n59) );
  AND2_X1 U137 ( .A1(n170), .A2(n91), .ZN(SUM[0]) );
  OR2_X1 U138 ( .A1(B[0]), .A2(A[0]), .ZN(n170) );
  OR2_X1 U139 ( .A1(A[11]), .A2(B[11]), .ZN(n171) );
  XNOR2_X1 U140 ( .A(n1), .B(n172), .ZN(SUM[11]) );
  AND2_X1 U141 ( .A1(n171), .A2(n43), .ZN(n172) );
  INV_X1 U142 ( .A(n98), .ZN(n173) );
  AND2_X1 U143 ( .A1(B[8]), .A2(A[8]), .ZN(n174) );
  INV_X1 U144 ( .A(n50), .ZN(n98) );
  OR2_X2 U145 ( .A1(A[8]), .A2(B[8]), .ZN(n186) );
  CLKBUF_X1 U146 ( .A(n43), .Z(n175) );
  NOR2_X1 U147 ( .A1(B[10]), .A2(A[10]), .ZN(n176) );
  NOR2_X1 U148 ( .A1(B[10]), .A2(A[10]), .ZN(n47) );
  OAI21_X1 U149 ( .B1(n51), .B2(n176), .A(n48), .ZN(n177) );
  AOI21_X1 U150 ( .B1(n45), .B2(n164), .A(n177), .ZN(n178) );
  AOI21_X1 U151 ( .B1(n45), .B2(n164), .A(n177), .ZN(n1) );
  XOR2_X1 U152 ( .A(n179), .B(n71), .Z(SUM[6]) );
  AND2_X1 U153 ( .A1(n181), .A2(n70), .ZN(n179) );
  XOR2_X1 U154 ( .A(n49), .B(n180), .Z(SUM[10]) );
  AND2_X1 U155 ( .A1(n97), .A2(n48), .ZN(n180) );
  OR2_X1 U156 ( .A1(B[6]), .A2(A[6]), .ZN(n181) );
  XNOR2_X1 U157 ( .A(n52), .B(n182), .ZN(SUM[9]) );
  AND2_X1 U158 ( .A1(n98), .A2(n51), .ZN(n182) );
  INV_X1 U159 ( .A(n38), .ZN(n36) );
  XNOR2_X1 U160 ( .A(n10), .B(n65), .ZN(SUM[7]) );
  INV_X1 U161 ( .A(n70), .ZN(n68) );
  OAI21_X1 U162 ( .B1(n43), .B2(n39), .A(n40), .ZN(n38) );
  OAI21_X1 U163 ( .B1(n74), .B2(n72), .A(n73), .ZN(n71) );
  NOR2_X1 U164 ( .A1(n42), .A2(n168), .ZN(n37) );
  XOR2_X1 U165 ( .A(n12), .B(n74), .Z(SUM[5]) );
  NAND2_X1 U166 ( .A1(n102), .A2(n73), .ZN(n12) );
  INV_X1 U167 ( .A(n72), .ZN(n102) );
  XOR2_X1 U168 ( .A(n60), .B(n9), .Z(SUM[8]) );
  INV_X1 U169 ( .A(n33), .ZN(n31) );
  NAND2_X1 U170 ( .A1(n95), .A2(n40), .ZN(n5) );
  NAND2_X1 U171 ( .A1(n183), .A2(n19), .ZN(n2) );
  NAND2_X1 U172 ( .A1(B[15]), .A2(A[15]), .ZN(n19) );
  NAND2_X1 U173 ( .A1(n166), .A2(n33), .ZN(n4) );
  XNOR2_X1 U174 ( .A(n27), .B(n3), .ZN(SUM[14]) );
  NAND2_X1 U175 ( .A1(n93), .A2(n26), .ZN(n3) );
  OR2_X1 U176 ( .A1(B[15]), .A2(A[15]), .ZN(n183) );
  AOI21_X1 U177 ( .B1(n187), .B2(n79), .A(n76), .ZN(n74) );
  INV_X1 U178 ( .A(n78), .ZN(n76) );
  OR2_X1 U179 ( .A1(B[7]), .A2(A[7]), .ZN(n184) );
  XOR2_X1 U180 ( .A(n14), .B(n82), .Z(SUM[3]) );
  NAND2_X1 U181 ( .A1(n104), .A2(n81), .ZN(n14) );
  INV_X1 U182 ( .A(n80), .ZN(n104) );
  OAI21_X1 U183 ( .B1(n80), .B2(n82), .A(n81), .ZN(n79) );
  NAND2_X1 U184 ( .A1(B[6]), .A2(A[6]), .ZN(n70) );
  NOR2_X1 U185 ( .A1(A[11]), .A2(B[11]), .ZN(n42) );
  OR2_X1 U186 ( .A1(B[2]), .A2(A[2]), .ZN(n185) );
  NOR2_X1 U187 ( .A1(B[5]), .A2(A[5]), .ZN(n72) );
  NAND2_X1 U188 ( .A1(A[13]), .A2(B[13]), .ZN(n33) );
  NOR2_X1 U189 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND2_X1 U190 ( .A1(B[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U191 ( .A1(B[5]), .A2(A[5]), .ZN(n73) );
  NAND2_X1 U192 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  NAND2_X1 U193 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  XNOR2_X1 U194 ( .A(n13), .B(n79), .ZN(SUM[4]) );
  NAND2_X1 U195 ( .A1(n187), .A2(n78), .ZN(n13) );
  NOR2_X1 U196 ( .A1(B[3]), .A2(A[3]), .ZN(n80) );
  AOI21_X1 U197 ( .B1(n87), .B2(n185), .A(n84), .ZN(n82) );
  INV_X1 U198 ( .A(n86), .ZN(n84) );
  NAND2_X1 U199 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  OR2_X1 U200 ( .A1(B[4]), .A2(A[4]), .ZN(n187) );
  XNOR2_X1 U201 ( .A(n15), .B(n87), .ZN(SUM[2]) );
  NAND2_X1 U202 ( .A1(n185), .A2(n86), .ZN(n15) );
  OAI21_X1 U203 ( .B1(n88), .B2(n91), .A(n89), .ZN(n87) );
  NOR2_X1 U204 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  NAND2_X1 U205 ( .A1(B[1]), .A2(A[1]), .ZN(n89) );
  XOR2_X1 U206 ( .A(n16), .B(n91), .Z(SUM[1]) );
  NAND2_X1 U207 ( .A1(n106), .A2(n89), .ZN(n16) );
  INV_X1 U208 ( .A(n88), .ZN(n106) );
  NAND2_X1 U209 ( .A1(B[0]), .A2(A[0]), .ZN(n91) );
  XNOR2_X1 U210 ( .A(n41), .B(n5), .ZN(SUM[12]) );
  AOI21_X1 U211 ( .B1(n38), .B2(n23), .A(n24), .ZN(n22) );
  NAND2_X1 U212 ( .A1(n37), .A2(n23), .ZN(n21) );
  NOR2_X1 U213 ( .A1(n32), .A2(n25), .ZN(n23) );
  INV_X1 U214 ( .A(n66), .ZN(n65) );
  AOI21_X1 U215 ( .B1(n181), .B2(n71), .A(n68), .ZN(n66) );
  NOR2_X1 U216 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  INV_X1 U217 ( .A(n25), .ZN(n93) );
  OAI21_X1 U218 ( .B1(n25), .B2(n33), .A(n26), .ZN(n24) );
  INV_X1 U219 ( .A(n168), .ZN(n95) );
  NAND2_X1 U220 ( .A1(B[3]), .A2(A[3]), .ZN(n81) );
  AOI21_X1 U221 ( .B1(n65), .B2(n184), .A(n62), .ZN(n60) );
  NAND2_X1 U222 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  NOR2_X1 U223 ( .A1(A[9]), .A2(B[9]), .ZN(n50) );
  XNOR2_X1 U224 ( .A(n20), .B(n2), .ZN(SUM[15]) );
  NAND2_X1 U225 ( .A1(B[14]), .A2(A[14]), .ZN(n26) );
  OAI21_X1 U226 ( .B1(n52), .B2(n173), .A(n51), .ZN(n49) );
  XNOR2_X1 U227 ( .A(n34), .B(n4), .ZN(SUM[13]) );
  INV_X1 U228 ( .A(n64), .ZN(n62) );
  NAND2_X1 U229 ( .A1(n184), .A2(n64), .ZN(n10) );
  NAND2_X1 U230 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  INV_X1 U231 ( .A(n53), .ZN(n52) );
  NAND2_X1 U232 ( .A1(n37), .A2(n166), .ZN(n28) );
  AOI21_X1 U233 ( .B1(n38), .B2(n166), .A(n31), .ZN(n29) );
  INV_X1 U234 ( .A(n163), .ZN(n97) );
  NOR2_X1 U235 ( .A1(n47), .A2(n50), .ZN(n45) );
  NAND2_X1 U236 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  OAI21_X1 U237 ( .B1(n167), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U238 ( .B1(n1), .B2(n28), .A(n29), .ZN(n27) );
  OAI21_X1 U239 ( .B1(n178), .B2(n42), .A(n175), .ZN(n41) );
  OAI21_X1 U240 ( .B1(n178), .B2(n165), .A(n36), .ZN(n34) );
  NAND2_X1 U241 ( .A1(n186), .A2(n59), .ZN(n9) );
  AOI21_X1 U242 ( .B1(n186), .B2(n62), .A(n174), .ZN(n55) );
  NAND2_X1 U243 ( .A1(n186), .A2(n184), .ZN(n54) );
endmodule


module recursive_add_layer_INPUT_SCALE4_WIDTH16_1 ( .in({\in[3][15] , 
        \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , \in[3][10] , 
        \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , \in[3][5] , \in[3][4] , 
        \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] , \in[2][15] , 
        \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , \in[2][10] , 
        \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , \in[2][5] , \in[2][4] , 
        \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] , \in[1][15] , 
        \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , \in[1][10] , 
        \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , 
        \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , 
        \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , 
        \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] , 
        \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), out );
  output [15:0] out;
  input \in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] ,
         \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] ,
         \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] ,
         \in[3][0] , \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] ,
         \in[2][11] , \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] ,
         \in[2][6] , \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] ,
         \in[2][1] , \in[2][0] , \in[1][15] , \in[1][14] , \in[1][13] ,
         \in[1][12] , \in[1][11] , \in[1][10] , \in[1][9] , \in[1][8] ,
         \in[1][7] , \in[1][6] , \in[1][5] , \in[1][4] , \in[1][3] ,
         \in[1][2] , \in[1][1] , \in[1][0] , \in[0][15] , \in[0][14] ,
         \in[0][13] , \in[0][12] , \in[0][11] , \in[0][10] , \in[0][9] ,
         \in[0][8] , \in[0][7] , \in[0][6] , \in[0][5] , \in[0][4] ,
         \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] ;
  wire   \genblk1.inter[1][15] , \genblk1.inter[1][14] ,
         \genblk1.inter[1][13] , \genblk1.inter[1][12] ,
         \genblk1.inter[1][11] , \genblk1.inter[1][10] , \genblk1.inter[1][9] ,
         \genblk1.inter[1][8] , \genblk1.inter[1][7] , \genblk1.inter[1][6] ,
         \genblk1.inter[1][5] , \genblk1.inter[1][4] , \genblk1.inter[1][3] ,
         \genblk1.inter[1][2] , \genblk1.inter[1][1] , \genblk1.inter[1][0] ,
         \genblk1.inter[0][15] , \genblk1.inter[0][14] ,
         \genblk1.inter[0][13] , \genblk1.inter[0][12] ,
         \genblk1.inter[0][11] , \genblk1.inter[0][10] , \genblk1.inter[0][9] ,
         \genblk1.inter[0][8] , \genblk1.inter[0][7] , \genblk1.inter[0][6] ,
         \genblk1.inter[0][5] , \genblk1.inter[0][4] , \genblk1.inter[0][3] ,
         \genblk1.inter[0][2] , \genblk1.inter[0][1] , \genblk1.inter[0][0] ;

  recursive_add_layer_INPUT_SCALE2_WIDTH16_1 \genblk1.next_layer  ( .in({
        \genblk1.inter[1][15] , \genblk1.inter[1][14] , \genblk1.inter[1][13] , 
        \genblk1.inter[1][12] , \genblk1.inter[1][11] , \genblk1.inter[1][10] , 
        \genblk1.inter[1][9] , \genblk1.inter[1][8] , \genblk1.inter[1][7] , 
        \genblk1.inter[1][6] , \genblk1.inter[1][5] , \genblk1.inter[1][4] , 
        \genblk1.inter[1][3] , \genblk1.inter[1][2] , \genblk1.inter[1][1] , 
        \genblk1.inter[1][0] , \genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }), .out(out) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_1_DW01_add_4 add_64_G2 ( .A({
        \in[2][15] , \in[2][14] , \in[2][13] , \in[2][12] , \in[2][11] , 
        \in[2][10] , \in[2][9] , \in[2][8] , \in[2][7] , \in[2][6] , 
        \in[2][5] , \in[2][4] , \in[2][3] , \in[2][2] , \in[2][1] , \in[2][0] }), .B({\in[3][15] , \in[3][14] , \in[3][13] , \in[3][12] , \in[3][11] , 
        \in[3][10] , \in[3][9] , \in[3][8] , \in[3][7] , \in[3][6] , 
        \in[3][5] , \in[3][4] , \in[3][3] , \in[3][2] , \in[3][1] , \in[3][0] }), .CI(1'b0), .SUM({\genblk1.inter[1][15] , \genblk1.inter[1][14] , 
        \genblk1.inter[1][13] , \genblk1.inter[1][12] , \genblk1.inter[1][11] , 
        \genblk1.inter[1][10] , \genblk1.inter[1][9] , \genblk1.inter[1][8] , 
        \genblk1.inter[1][7] , \genblk1.inter[1][6] , \genblk1.inter[1][5] , 
        \genblk1.inter[1][4] , \genblk1.inter[1][3] , \genblk1.inter[1][2] , 
        \genblk1.inter[1][1] , \genblk1.inter[1][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_1_DW01_add_5 add_64 ( .A({
        \in[0][15] , \in[0][14] , \in[0][13] , \in[0][12] , \in[0][11] , 
        \in[0][10] , \in[0][9] , \in[0][8] , \in[0][7] , \in[0][6] , 
        \in[0][5] , \in[0][4] , \in[0][3] , \in[0][2] , \in[0][1] , \in[0][0] }), .B({\in[1][15] , \in[1][14] , \in[1][13] , \in[1][12] , \in[1][11] , 
        \in[1][10] , \in[1][9] , \in[1][8] , \in[1][7] , \in[1][6] , 
        \in[1][5] , \in[1][4] , \in[1][3] , \in[1][2] , \in[1][1] , \in[1][0] }), .CI(1'b0), .SUM({\genblk1.inter[0][15] , \genblk1.inter[0][14] , 
        \genblk1.inter[0][13] , \genblk1.inter[0][12] , \genblk1.inter[0][11] , 
        \genblk1.inter[0][10] , \genblk1.inter[0][9] , \genblk1.inter[0][8] , 
        \genblk1.inter[0][7] , \genblk1.inter[0][6] , \genblk1.inter[0][5] , 
        \genblk1.inter[0][4] , \genblk1.inter[0][3] , \genblk1.inter[0][2] , 
        \genblk1.inter[0][1] , \genblk1.inter[0][0] }) );
endmodule


module element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_1 ( .a({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , 
        \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , 
        \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .x({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , 
        \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] , \x[2][5] , 
        \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , \x[1][7] , 
        \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , 
        \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , 
        \x[0][2] , \x[0][1] , \x[0][0] }), y );
  output [15:0] y;
  input \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] ,
         \a[3][1] , \a[3][0] , \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] ,
         \a[2][3] , \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] ,
         \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] ,
         \a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] ,
         \a[0][1] , \a[0][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , \x[2][6] ,
         \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] ,
         \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] ,
         \x[1][1] , \x[1][0] , \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] ;
  wire   \multout[3][15] , \multout[3][14] , \multout[3][13] ,
         \multout[3][12] , \multout[3][11] , \multout[3][10] , \multout[3][9] ,
         \multout[3][8] , \multout[3][7] , \multout[3][6] , \multout[3][5] ,
         \multout[3][4] , \multout[3][3] , \multout[3][2] , \multout[3][1] ,
         \multout[3][0] , \multout[2][15] , \multout[2][14] , \multout[2][13] ,
         \multout[2][12] , \multout[2][11] , \multout[2][10] , \multout[2][9] ,
         \multout[2][8] , \multout[2][7] , \multout[2][6] , \multout[2][5] ,
         \multout[2][4] , \multout[2][3] , \multout[2][2] , \multout[2][1] ,
         \multout[2][0] , \multout[1][15] , \multout[1][14] , \multout[1][13] ,
         \multout[1][12] , \multout[1][11] , \multout[1][10] , \multout[1][9] ,
         \multout[1][8] , \multout[1][7] , \multout[1][6] , \multout[1][5] ,
         \multout[1][4] , \multout[1][3] , \multout[1][2] , \multout[1][1] ,
         \multout[1][0] , \multout[0][15] , \multout[0][14] , \multout[0][13] ,
         \multout[0][12] , \multout[0][11] , \multout[0][10] , \multout[0][9] ,
         \multout[0][8] , \multout[0][7] , \multout[0][6] , \multout[0][5] ,
         \multout[0][4] , \multout[0][3] , \multout[0][2] , \multout[0][1] ,
         \multout[0][0] ;

  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_4 \genblk1[0].mult  ( .ia({\a[0][7] , 
        \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , 
        \a[0][0] }), .ix({\x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , 
        \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] }), .out({\multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_3 \genblk1[1].mult  ( .ia({\a[1][7] , 
        \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , 
        \a[1][0] }), .ix({\x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , 
        \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] }), .out({\multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_2 \genblk1[2].mult  ( .ia({\a[2][7] , 
        \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , \a[2][1] , 
        \a[2][0] }), .ix({\x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] , 
        \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] }), .out({\multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] }) );
  mult_layer_INPUT_WIDTH8_OUTPUT_WIDTH16_1 \genblk1[3].mult  ( .ia({\a[3][7] , 
        \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , 
        \a[3][0] }), .ix({\x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] , 
        \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] }), .out({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] }) );
  recursive_add_layer_INPUT_SCALE4_WIDTH16_1 add ( .in({\multout[3][15] , 
        \multout[3][14] , \multout[3][13] , \multout[3][12] , \multout[3][11] , 
        \multout[3][10] , \multout[3][9] , \multout[3][8] , \multout[3][7] , 
        \multout[3][6] , \multout[3][5] , \multout[3][4] , \multout[3][3] , 
        \multout[3][2] , \multout[3][1] , \multout[3][0] , \multout[2][15] , 
        \multout[2][14] , \multout[2][13] , \multout[2][12] , \multout[2][11] , 
        \multout[2][10] , \multout[2][9] , \multout[2][8] , \multout[2][7] , 
        \multout[2][6] , \multout[2][5] , \multout[2][4] , \multout[2][3] , 
        \multout[2][2] , \multout[2][1] , \multout[2][0] , \multout[1][15] , 
        \multout[1][14] , \multout[1][13] , \multout[1][12] , \multout[1][11] , 
        \multout[1][10] , \multout[1][9] , \multout[1][8] , \multout[1][7] , 
        \multout[1][6] , \multout[1][5] , \multout[1][4] , \multout[1][3] , 
        \multout[1][2] , \multout[1][1] , \multout[1][0] , \multout[0][15] , 
        \multout[0][14] , \multout[0][13] , \multout[0][12] , \multout[0][11] , 
        \multout[0][10] , \multout[0][9] , \multout[0][8] , \multout[0][7] , 
        \multout[0][6] , \multout[0][5] , \multout[0][4] , \multout[0][3] , 
        \multout[0][2] , \multout[0][1] , \multout[0][0] }), .out(y) );
endmodule


module data_path_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16 ( clk, en_a, en_x, 
        en_y, clr_addr_a, clr_addr_x, clr_addr_y, of_a, of_x, of_y, data_in, 
        data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y;
  output of_a, of_x, of_y;
  wire   N22, N23, \a[15][7] , \a[15][6] , \a[15][5] , \a[15][4] , \a[15][2] ,
         \a[15][1] , \a[15][0] , \a[14][7] , \a[14][6] , \a[14][5] ,
         \a[14][4] , \a[14][3] , \a[14][2] , \a[14][1] , \a[14][0] ,
         \a[13][6] , \a[13][5] , \a[13][4] , \a[13][3] , \a[13][2] ,
         \a[13][1] , \a[13][0] , \a[12][6] , \a[12][5] , \a[12][4] ,
         \a[12][3] , \a[12][2] , \a[12][1] , \a[12][0] , \a[11][7] ,
         \a[11][6] , \a[11][5] , \a[11][4] , \a[11][3] , \a[11][2] ,
         \a[11][1] , \a[11][0] , \a[10][6] , \a[10][5] , \a[10][4] ,
         \a[10][2] , \a[10][1] , \a[10][0] , \a[9][6] , \a[9][5] , \a[9][4] ,
         \a[9][3] , \a[9][2] , \a[9][1] , \a[9][0] , \a[8][7] , \a[8][6] ,
         \a[8][5] , \a[8][4] , \a[8][3] , \a[8][2] , \a[8][1] , \a[8][0] ,
         \a[7][6] , \a[7][5] , \a[7][4] , \a[7][3] , \a[7][2] , \a[7][0] ,
         \a[6][7] , \a[6][6] , \a[6][5] , \a[6][4] , \a[6][3] , \a[6][2] ,
         \a[6][1] , \a[6][0] , \a[5][7] , \a[5][6] , \a[5][5] , \a[5][4] ,
         \a[5][2] , \a[5][1] , \a[5][0] , \a[4][7] , \a[4][6] , \a[4][5] ,
         \a[4][4] , \a[4][2] , \a[4][1] , \a[4][0] , \a[3][7] , \a[3][6] ,
         \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , \a[3][1] , \a[3][0] ,
         \a[2][7] , \a[2][6] , \a[2][5] , \a[2][4] , \a[2][2] , \a[2][1] ,
         \a[2][0] , \a[1][7] , \a[1][6] , \a[1][5] , \a[1][4] , \a[1][3] ,
         \a[1][2] , \a[1][1] , \a[1][0] , \a[0][7] , \a[0][6] , \a[0][5] ,
         \a[0][4] , \a[0][3] , \a[0][2] , \a[0][1] , \a[0][0] , \x[3][7] ,
         \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] ,
         \x[3][0] , \x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] , \x[2][3] ,
         \x[2][2] , \x[2][1] , \x[2][0] , \x[1][7] , \x[1][6] , \x[1][5] ,
         \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] , \x[0][7] ,
         \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] ,
         \x[0][0] , \y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] , \y[3][11] ,
         \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] , \y[3][5] ,
         \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] , \y[2][15] ,
         \y[2][14] , \y[2][13] , \y[2][12] , \y[2][11] , \y[2][10] , \y[2][9] ,
         \y[2][8] , \y[2][7] , \y[2][6] , \y[2][5] , \y[2][4] , \y[2][3] ,
         \y[2][2] , \y[2][1] , \y[2][0] , \y[1][15] , \y[1][14] , \y[1][13] ,
         \y[1][12] , \y[1][11] , \y[1][10] , \y[1][9] , \y[1][8] , \y[1][7] ,
         \y[1][6] , \y[1][5] , \y[1][4] , \y[1][3] , \y[1][2] , \y[1][1] ,
         \y[1][0] , \y[0][15] , \y[0][14] , \y[0][13] , \y[0][12] , \y[0][11] ,
         \y[0][10] , \y[0][9] , \y[0][8] , \y[0][7] , \y[0][6] , \y[0][5] ,
         \y[0][4] , \y[0][3] , \y[0][2] , \y[0][1] , \y[0][0] , N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N79, N80, N81, N87, N89,
         N90, N94, N95, N99, N100, N103, N104, N105, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n12, n15, n16, n40, n50, n60, n70, n71, n81, n109,
         n119, n193, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n11, n13, n14, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429;
  wire   [3:0] addr_a;
  wire   [1:0] addr_x;
  assign of_a = N103;
  assign of_x = N104;
  assign of_y = N105;

  DFF_X1 \data_out_reg[15]  ( .D(N66), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N67), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N68), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N69), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N70), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N71), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N72), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N73), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N74), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N75), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N76), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N77), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N79), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N80), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N81), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \addr_a_reg[0]  ( .D(N87), .CK(clk), .Q(addr_a[0]) );
  DFF_X1 \a_reg[3][6]  ( .D(n344), .CK(clk), .Q(\a[3][6] ) );
  DFF_X1 \a_reg[3][4]  ( .D(n346), .CK(clk), .Q(\a[3][4] ) );
  DFF_X1 \a_reg[3][2]  ( .D(n348), .CK(clk), .Q(\a[3][2] ) );
  DFF_X1 \a_reg[3][0]  ( .D(n350), .CK(clk), .Q(\a[3][0] ) );
  DFF_X1 \a_reg[2][6]  ( .D(n352), .CK(clk), .Q(\a[2][6] ) );
  DFF_X1 \a_reg[2][4]  ( .D(n354), .CK(clk), .Q(\a[2][4] ) );
  DFF_X1 \a_reg[2][2]  ( .D(n356), .CK(clk), .Q(\a[2][2] ), .QN(n52) );
  DFF_X1 \a_reg[2][0]  ( .D(n358), .CK(clk), .Q(\a[2][0] ) );
  DFF_X1 \a_reg[1][6]  ( .D(n360), .CK(clk), .Q(\a[1][6] ) );
  DFF_X1 \a_reg[1][4]  ( .D(n362), .CK(clk), .Q(\a[1][4] ) );
  DFF_X1 \a_reg[1][2]  ( .D(n364), .CK(clk), .Q(\a[1][2] ) );
  DFF_X1 \a_reg[1][0]  ( .D(n366), .CK(clk), .Q(\a[1][0] ) );
  DFF_X1 \a_reg[0][6]  ( .D(n368), .CK(clk), .Q(\a[0][6] ) );
  DFF_X1 \a_reg[0][4]  ( .D(n370), .CK(clk), .Q(\a[0][4] ), .QN(n106) );
  DFF_X1 \a_reg[0][2]  ( .D(n372), .CK(clk), .Q(\a[0][2] ) );
  DFF_X1 \a_reg[0][0]  ( .D(n374), .CK(clk), .Q(\a[0][0] ) );
  DFF_X1 \a_reg[11][6]  ( .D(n280), .CK(clk), .Q(\a[11][6] ) );
  DFF_X1 \a_reg[11][4]  ( .D(n282), .CK(clk), .Q(\a[11][4] ) );
  DFF_X1 \a_reg[11][2]  ( .D(n284), .CK(clk), .Q(\a[11][2] ) );
  DFF_X1 \a_reg[11][0]  ( .D(n286), .CK(clk), .Q(\a[11][0] ) );
  DFF_X1 \a_reg[10][7]  ( .D(n287), .CK(clk), .QN(n144) );
  DFF_X1 \a_reg[10][6]  ( .D(n288), .CK(clk), .Q(\a[10][6] ) );
  DFF_X1 \a_reg[10][4]  ( .D(n290), .CK(clk), .Q(\a[10][4] ) );
  DFF_X1 \a_reg[10][2]  ( .D(n292), .CK(clk), .Q(\a[10][2] ) );
  DFF_X1 \a_reg[10][0]  ( .D(n294), .CK(clk), .Q(\a[10][0] ) );
  DFF_X1 \a_reg[9][6]  ( .D(n296), .CK(clk), .Q(\a[9][6] ) );
  DFF_X1 \a_reg[9][4]  ( .D(n298), .CK(clk), .Q(\a[9][4] ) );
  DFF_X1 \a_reg[9][2]  ( .D(n300), .CK(clk), .Q(\a[9][2] ) );
  DFF_X1 \a_reg[9][0]  ( .D(n302), .CK(clk), .Q(\a[9][0] ) );
  DFF_X1 \a_reg[8][6]  ( .D(n304), .CK(clk), .Q(\a[8][6] ) );
  DFF_X1 \a_reg[8][4]  ( .D(n306), .CK(clk), .Q(\a[8][4] ) );
  DFF_X1 \a_reg[8][2]  ( .D(n308), .CK(clk), .Q(\a[8][2] ) );
  DFF_X1 \a_reg[8][0]  ( .D(n310), .CK(clk), .Q(\a[8][0] ) );
  DFF_X1 \a_reg[7][6]  ( .D(n312), .CK(clk), .Q(\a[7][6] ) );
  DFF_X1 \a_reg[7][4]  ( .D(n314), .CK(clk), .Q(\a[7][4] ) );
  DFF_X1 \a_reg[7][2]  ( .D(n316), .CK(clk), .Q(\a[7][2] ) );
  DFF_X1 \a_reg[7][0]  ( .D(n318), .CK(clk), .Q(\a[7][0] ) );
  DFF_X1 \a_reg[6][6]  ( .D(n320), .CK(clk), .Q(\a[6][6] ) );
  DFF_X1 \a_reg[6][4]  ( .D(n322), .CK(clk), .Q(\a[6][4] ) );
  DFF_X1 \a_reg[6][2]  ( .D(n324), .CK(clk), .Q(\a[6][2] ) );
  DFF_X1 \a_reg[6][0]  ( .D(n326), .CK(clk), .Q(\a[6][0] ) );
  DFF_X1 \a_reg[5][6]  ( .D(n328), .CK(clk), .Q(\a[5][6] ) );
  DFF_X1 \a_reg[5][4]  ( .D(n330), .CK(clk), .Q(\a[5][4] ) );
  DFF_X1 \a_reg[5][2]  ( .D(n332), .CK(clk), .Q(\a[5][2] ) );
  DFF_X1 \a_reg[5][0]  ( .D(n334), .CK(clk), .Q(\a[5][0] ) );
  DFF_X1 \a_reg[4][6]  ( .D(n336), .CK(clk), .Q(\a[4][6] ) );
  DFF_X1 \a_reg[4][4]  ( .D(n338), .CK(clk), .Q(\a[4][4] ) );
  DFF_X1 \a_reg[4][2]  ( .D(n340), .CK(clk), .Q(\a[4][2] ) );
  DFF_X1 \a_reg[4][0]  ( .D(n342), .CK(clk), .Q(\a[4][0] ) );
  DFF_X1 \a_reg[14][6]  ( .D(n256), .CK(clk), .Q(\a[14][6] ) );
  DFF_X1 \a_reg[14][5]  ( .D(n257), .CK(clk), .Q(\a[14][5] ), .QN(n54) );
  DFF_X1 \a_reg[14][4]  ( .D(n258), .CK(clk), .Q(\a[14][4] ) );
  DFF_X1 \a_reg[14][2]  ( .D(n260), .CK(clk), .Q(\a[14][2] ) );
  DFF_X1 \a_reg[14][0]  ( .D(n262), .CK(clk), .Q(\a[14][0] ) );
  DFF_X1 \a_reg[13][6]  ( .D(n264), .CK(clk), .Q(\a[13][6] ) );
  DFF_X1 \a_reg[13][4]  ( .D(n266), .CK(clk), .Q(\a[13][4] ) );
  DFF_X1 \a_reg[13][2]  ( .D(n268), .CK(clk), .Q(\a[13][2] ) );
  DFF_X1 \a_reg[13][0]  ( .D(n270), .CK(clk), .Q(\a[13][0] ) );
  DFF_X1 \a_reg[12][2]  ( .D(n276), .CK(clk), .Q(\a[12][2] ) );
  DFF_X1 \a_reg[12][0]  ( .D(n278), .CK(clk), .Q(\a[12][0] ) );
  DFF_X1 \a_reg[12][6]  ( .D(n272), .CK(clk), .Q(\a[12][6] ) );
  DFF_X1 \a_reg[12][4]  ( .D(n274), .CK(clk), .Q(\a[12][4] ) );
  DFF_X1 \a_reg[15][6]  ( .D(n248), .CK(clk), .Q(\a[15][6] ) );
  DFF_X1 \a_reg[15][4]  ( .D(n250), .CK(clk), .Q(\a[15][4] ) );
  DFF_X1 \a_reg[15][2]  ( .D(n252), .CK(clk), .Q(\a[15][2] ) );
  DFF_X1 \a_reg[15][0]  ( .D(n254), .CK(clk), .Q(\a[15][0] ) );
  DFF_X1 \x_reg[1][1]  ( .D(n237), .CK(clk), .Q(\x[1][1] ), .QN(n187) );
  DFF_X1 \x_reg[1][0]  ( .D(n238), .CK(clk), .Q(\x[1][0] ) );
  DFF_X1 \x_reg[0][6]  ( .D(n240), .CK(clk), .Q(\x[0][6] ), .QN(n169) );
  DFF_X1 \x_reg[0][5]  ( .D(n241), .CK(clk), .Q(\x[0][5] ), .QN(n177) );
  DFF_X1 \x_reg[0][0]  ( .D(n246), .CK(clk), .Q(\x[0][0] ) );
  DFF_X1 \x_reg[2][2]  ( .D(n228), .CK(clk), .Q(\x[2][2] ) );
  DFF_X1 \x_reg[2][1]  ( .D(n229), .CK(clk), .Q(\x[2][1] ), .QN(n30) );
  DFF_X1 \x_reg[2][0]  ( .D(n230), .CK(clk), .Q(\x[2][0] ), .QN(n99) );
  DFF_X1 \x_reg[3][6]  ( .D(n216), .CK(clk), .Q(\x[3][6] ), .QN(n2) );
  DFF_X1 \x_reg[3][5]  ( .D(n217), .CK(clk), .Q(\x[3][5] ), .QN(n3) );
  DFF_X1 \x_reg[3][0]  ( .D(n222), .CK(clk), .Q(\x[3][0] ), .QN(n8) );
  XOR2_X1 U373 ( .A(n15), .B(addr_x[0]), .Z(n207) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_0 \genblk1[0].element  ( 
        .a({n172, \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , \a[3][2] , 
        \a[3][1] , \a[3][0] , n161, \a[2][6] , n199, \a[2][4] , n186, 
        \a[2][2] , \a[2][1] , \a[2][0] , \a[1][7] , \a[1][6] , n103, \a[1][4] , 
        n88, \a[1][2] , n84, \a[1][0] , n90, \a[0][6] , n147, \a[0][4] , 
        \a[0][3] , \a[0][2] , n184, \a[0][0] }), .x({n32, n404, n407, 
        \x[3][4] , \x[3][3] , \x[3][2] , n74, \x[3][0] , \x[2][7] , \x[2][6] , 
        \x[2][5] , \x[2][4] , \x[2][3] , n405, n31, \x[2][0] , \x[1][7] , 
        \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , n188, n408, 
        \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , \x[0][2] , 
        \x[0][1] , \x[0][0] }), .y({\y[0][15] , \y[0][14] , \y[0][13] , 
        \y[0][12] , \y[0][11] , \y[0][10] , \y[0][9] , \y[0][8] , \y[0][7] , 
        \y[0][6] , \y[0][5] , \y[0][4] , \y[0][3] , \y[0][2] , \y[0][1] , 
        \y[0][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_3 \genblk1[1].element  ( 
        .a({n165, \a[7][6] , \a[7][5] , \a[7][4] , n190, \a[7][2] , n105, 
        \a[7][0] , n51, \a[6][6] , \a[6][5] , \a[6][4] , \a[6][3] , \a[6][2] , 
        \a[6][1] , \a[6][0] , \a[5][7] , \a[5][6] , n157, \a[5][4] , n92, 
        \a[5][2] , n201, \a[5][0] , n167, \a[4][6] , n163, \a[4][4] , n203, 
        \a[4][2] , n69, \a[4][0] }), .x({\x[3][7] , n404, n407, \x[3][4] , n42, 
        \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , n38, n44, n65, n61, n405, 
        n31, n100, \x[1][7] , n46, n48, \x[1][4] , \x[1][3] , \x[1][2] , 
        \x[1][1] , \x[1][0] , n21, \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , 
        \x[0][2] , \x[0][1] , \x[0][0] }), .y({\y[1][15] , \y[1][14] , 
        \y[1][13] , \y[1][12] , \y[1][11] , \y[1][10] , \y[1][9] , \y[1][8] , 
        \y[1][7] , \y[1][6] , \y[1][5] , \y[1][4] , \y[1][3] , \y[1][2] , 
        \y[1][1] , \y[1][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_2 \genblk1[2].element  ( 
        .a({n17, \a[11][6] , \a[11][5] , \a[11][4] , \a[11][3] , \a[11][2] , 
        n197, \a[11][0] , n145, \a[10][6] , \a[10][5] , \a[10][4] , n135, 
        \a[10][2] , \a[10][1] , \a[10][0] , n139, \a[9][6] , n143, \a[9][4] , 
        n155, \a[9][2] , \a[9][1] , \a[9][0] , \a[8][7] , \a[8][6] , n149, 
        \a[8][4] , \a[8][3] , \a[8][2] , \a[8][1] , \a[8][0] }), .x({n32, n72, 
        n73, \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , 
        n38, n44, n65, n61, n405, n406, n100, \x[1][7] , \x[1][6] , \x[1][5] , 
        \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , n408, \x[0][7] , n170, 
        n178, \x[0][4] , \x[0][3] , \x[0][2] , n23, \x[0][0] }), .y({
        \y[2][15] , \y[2][14] , \y[2][13] , \y[2][12] , \y[2][11] , \y[2][10] , 
        \y[2][9] , \y[2][8] , \y[2][7] , \y[2][6] , \y[2][5] , \y[2][4] , 
        \y[2][3] , \y[2][2] , \y[2][1] , \y[2][0] }) );
  element_layer_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16_1 \genblk1[3].element  ( 
        .a({n159, \a[15][6] , n141, \a[15][4] , n137, \a[15][2] , n153, 
        \a[15][0] , \a[14][7] , \a[14][6] , \a[14][5] , \a[14][4] , n63, 
        \a[14][2] , \a[14][1] , \a[14][0] , n82, \a[13][6] , n78, \a[13][4] , 
        n174, \a[13][2] , \a[13][1] , \a[13][0] , n95, \a[12][6] , n76, 
        \a[12][4] , n192, \a[12][2] , n151, \a[12][0] }), .x({\x[3][7] , n72, 
        n73, \x[3][4] , n42, \x[3][2] , \x[3][1] , \x[3][0] , \x[2][7] , 
        \x[2][6] , \x[2][5] , \x[2][4] , \x[2][3] , n405, n406, \x[2][0] , 
        \x[1][7] , n46, n48, \x[1][4] , \x[1][3] , \x[1][2] , n188, \x[1][0] , 
        n21, n170, n178, \x[0][4] , \x[0][3] , \x[0][2] , n23, \x[0][0] }), 
        .y({\y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] , \y[3][11] , 
        \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] , \y[3][5] , 
        \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] }) );
  DFF_X2 \a_reg[8][7]  ( .D(n303), .CK(clk), .Q(\a[8][7] ) );
  DFF_X2 \x_reg[3][1]  ( .D(n221), .CK(clk), .Q(\x[3][1] ), .QN(n7) );
  DFF_X1 \a_reg[0][3]  ( .D(n371), .CK(clk), .Q(\a[0][3] ), .QN(n175) );
  DFF_X1 \a_reg[3][3]  ( .D(n347), .CK(clk), .Q(\a[3][3] ), .QN(n181) );
  DFF_X1 \a_reg[6][3]  ( .D(n323), .CK(clk), .Q(\a[6][3] ), .QN(n179) );
  DFF_X1 \a_reg[10][1]  ( .D(n293), .CK(clk), .Q(\a[10][1] ), .QN(n18) );
  DFF_X2 \a_reg[7][5]  ( .D(n313), .CK(clk), .Q(\a[7][5] ), .QN(n194) );
  DFF_X1 \a_reg[6][1]  ( .D(n325), .CK(clk), .Q(\a[6][1] ) );
  DFF_X1 \a_reg[4][3]  ( .D(n339), .CK(clk), .QN(n202) );
  DFF_X1 \a_reg[8][3]  ( .D(n307), .CK(clk), .Q(\a[8][3] ) );
  DFF_X1 \a_reg[3][1]  ( .D(n349), .CK(clk), .Q(\a[3][1] ), .QN(n57) );
  DFF_X1 \a_reg[5][1]  ( .D(n333), .CK(clk), .Q(\a[5][1] ), .QN(n200) );
  DFF_X1 \a_reg[2][1]  ( .D(n357), .CK(clk), .Q(\a[2][1] ), .QN(n33) );
  DFF_X1 \a_reg[2][5]  ( .D(n353), .CK(clk), .Q(\a[2][5] ), .QN(n198) );
  DFF_X1 \a_reg[11][1]  ( .D(n285), .CK(clk), .Q(\a[11][1] ), .QN(n196) );
  DFF_X1 \a_reg[14][1]  ( .D(n261), .CK(clk), .Q(\a[14][1] ), .QN(n28) );
  DFF_X1 \a_reg[12][3]  ( .D(n275), .CK(clk), .Q(\a[12][3] ), .QN(n191) );
  DFF_X1 \a_reg[7][3]  ( .D(n315), .CK(clk), .Q(\a[7][3] ), .QN(n189) );
  DFF_X1 \a_reg[8][1]  ( .D(n309), .CK(clk), .Q(\a[8][1] ) );
  DFF_X1 \a_reg[0][1]  ( .D(n373), .CK(clk), .Q(\a[0][1] ), .QN(n183) );
  DFF_X1 \a_reg[13][3]  ( .D(n267), .CK(clk), .Q(\a[13][3] ), .QN(n173) );
  DFF_X1 \a_reg[3][7]  ( .D(n343), .CK(clk), .Q(\a[3][7] ), .QN(n171) );
  DFF_X1 \a_reg[9][1]  ( .D(n301), .CK(clk), .Q(\a[9][1] ), .QN(n11) );
  DFF_X2 \x_reg[3][2]  ( .D(n220), .CK(clk), .Q(\x[3][2] ), .QN(n6) );
  DFF_X1 \a_reg[13][7]  ( .D(n263), .CK(clk), .Q(n82) );
  DFF_X1 \a_reg[4][7]  ( .D(n335), .CK(clk), .Q(\a[4][7] ), .QN(n166) );
  DFF_X2 \x_reg[3][4]  ( .D(n218), .CK(clk), .Q(\x[3][4] ), .QN(n4) );
  DFF_X1 \a_reg[7][7]  ( .D(n311), .CK(clk), .QN(n164) );
  DFF_X1 \a_reg[13][1]  ( .D(n269), .CK(clk), .Q(\a[13][1] ), .QN(n24) );
  DFF_X2 \x_reg[1][3]  ( .D(n235), .CK(clk), .Q(\x[1][3] ) );
  DFF_X1 \a_reg[4][5]  ( .D(n337), .CK(clk), .Q(\a[4][5] ), .QN(n162) );
  DFF_X2 \x_reg[0][3]  ( .D(n243), .CK(clk), .Q(\x[0][3] ) );
  DFF_X1 \a_reg[2][7]  ( .D(n351), .CK(clk), .Q(\a[2][7] ), .QN(n160) );
  DFF_X1 \a_reg[15][7]  ( .D(n247), .CK(clk), .Q(\a[15][7] ), .QN(n158) );
  DFF_X1 \a_reg[5][5]  ( .D(n329), .CK(clk), .Q(\a[5][5] ), .QN(n156) );
  DFF_X1 \a_reg[9][3]  ( .D(n299), .CK(clk), .Q(\a[9][3] ), .QN(n154) );
  DFF_X1 \a_reg[15][1]  ( .D(n253), .CK(clk), .Q(\a[15][1] ), .QN(n152) );
  DFF_X1 \a_reg[12][1]  ( .D(n277), .CK(clk), .Q(\a[12][1] ), .QN(n150) );
  DFF_X1 \a_reg[8][5]  ( .D(n305), .CK(clk), .Q(\a[8][5] ), .QN(n148) );
  DFF_X1 \a_reg[0][5]  ( .D(n369), .CK(clk), .Q(\a[0][5] ), .QN(n146) );
  DFF_X2 \x_reg[2][7]  ( .D(n223), .CK(clk), .Q(\x[2][7] ) );
  DFF_X1 \a_reg[9][5]  ( .D(n297), .CK(clk), .Q(\a[9][5] ), .QN(n142) );
  DFF_X1 \a_reg[15][5]  ( .D(n249), .CK(clk), .Q(\a[15][5] ), .QN(n140) );
  DFF_X1 \addr_y_reg[0]  ( .D(N99), .CK(clk), .Q(N22), .QN(n427) );
  DFF_X1 \addr_x_reg[0]  ( .D(N94), .CK(clk), .Q(addr_x[0]), .QN(n16) );
  DFF_X1 \addr_y_reg[1]  ( .D(N100), .CK(clk), .Q(N23), .QN(n426) );
  DFF_X1 \addr_x_reg[1]  ( .D(N95), .CK(clk), .Q(addr_x[1]), .QN(n15) );
  DFF_X1 \addr_a_reg[2]  ( .D(N89), .CK(clk), .Q(addr_a[2]), .QN(n10) );
  DFF_X1 \addr_a_reg[1]  ( .D(n428), .CK(clk), .Q(addr_a[1]), .QN(n12) );
  DFF_X1 \addr_a_reg[3]  ( .D(N90), .CK(clk), .Q(addr_a[3]), .QN(n9) );
  SDFF_X1 \data_out_reg[3]  ( .D(n379), .SI(n378), .SE(N23), .CK(clk), .Q(
        data_out[3]) );
  DFF_X1 \a_reg[9][7]  ( .D(n295), .CK(clk), .Q(n96), .QN(n138) );
  DFF_X1 \a_reg[3][5]  ( .D(n345), .CK(clk), .Q(\a[3][5] ), .QN(n39) );
  DFF_X2 \x_reg[0][2]  ( .D(n244), .CK(clk), .Q(\x[0][2] ) );
  DFF_X1 \a_reg[11][5]  ( .D(n281), .CK(clk), .Q(\a[11][5] ), .QN(n85) );
  DFF_X1 \a_reg[11][3]  ( .D(n283), .CK(clk), .Q(\a[11][3] ) );
  DFF_X1 \a_reg[14][7]  ( .D(n255), .CK(clk), .Q(\a[14][7] ), .QN(n35) );
  DFF_X2 \x_reg[0][4]  ( .D(n242), .CK(clk), .Q(\x[0][4] ) );
  DFF_X2 \x_reg[1][4]  ( .D(n234), .CK(clk), .Q(\x[1][4] ) );
  DFF_X1 \a_reg[15][3]  ( .D(n251), .CK(clk), .Q(n80), .QN(n136) );
  DFF_X1 \a_reg[10][3]  ( .D(n291), .CK(clk), .QN(n134) );
  DFF_X1 \a_reg[10][5]  ( .D(n289), .CK(clk), .Q(\a[10][5] ), .QN(n97) );
  DFF_X1 \a_reg[7][1]  ( .D(n317), .CK(clk), .QN(n104) );
  DFF_X1 \a_reg[1][5]  ( .D(n361), .CK(clk), .Q(\a[1][5] ), .QN(n102) );
  DFF_X2 \x_reg[1][7]  ( .D(n231), .CK(clk), .Q(\x[1][7] ) );
  DFF_X1 \a_reg[12][7]  ( .D(n271), .CK(clk), .QN(n94) );
  DFF_X1 \a_reg[5][3]  ( .D(n331), .CK(clk), .QN(n91) );
  DFF_X2 \x_reg[1][2]  ( .D(n236), .CK(clk), .Q(\x[1][2] ) );
  DFF_X1 \a_reg[0][7]  ( .D(n367), .CK(clk), .Q(\a[0][7] ), .QN(n89) );
  DFF_X1 \a_reg[1][3]  ( .D(n363), .CK(clk), .Q(\a[1][3] ), .QN(n87) );
  DFF_X1 \a_reg[1][1]  ( .D(n365), .CK(clk), .Q(\a[1][1] ), .QN(n83) );
  DFF_X2 \a_reg[1][7]  ( .D(n359), .CK(clk), .Q(\a[1][7] ) );
  DFF_X1 \a_reg[13][5]  ( .D(n265), .CK(clk), .Q(\a[13][5] ), .QN(n77) );
  DFF_X1 \a_reg[12][5]  ( .D(n273), .CK(clk), .Q(\a[12][5] ), .QN(n75) );
  DFF_X1 \a_reg[4][1]  ( .D(n341), .CK(clk), .Q(\a[4][1] ), .QN(n68) );
  DFF_X1 \a_reg[5][7]  ( .D(n327), .CK(clk), .Q(\a[5][7] ), .QN(n66) );
  DFF_X1 \x_reg[2][4]  ( .D(n226), .CK(clk), .Q(\x[2][4] ), .QN(n64) );
  DFF_X1 \a_reg[14][3]  ( .D(n259), .CK(clk), .Q(\a[14][3] ), .QN(n62) );
  DFF_X1 \x_reg[2][3]  ( .D(n227), .CK(clk), .Q(\x[2][3] ), .QN(n59) );
  DFF_X1 \a_reg[6][5]  ( .D(n321), .CK(clk), .Q(\a[6][5] ), .QN(n26) );
  DFF_X1 \a_reg[6][7]  ( .D(n319), .CK(clk), .Q(\a[6][7] ), .QN(n49) );
  DFF_X1 \x_reg[1][5]  ( .D(n233), .CK(clk), .Q(\x[1][5] ), .QN(n47) );
  DFF_X1 \x_reg[1][6]  ( .D(n232), .CK(clk), .Q(\x[1][6] ), .QN(n45) );
  DFF_X1 \x_reg[2][5]  ( .D(n225), .CK(clk), .Q(\x[2][5] ), .QN(n43) );
  DFF_X1 \x_reg[3][3]  ( .D(n219), .CK(clk), .Q(\x[3][3] ), .QN(n5) );
  DFF_X1 \x_reg[2][6]  ( .D(n224), .CK(clk), .Q(\x[2][6] ), .QN(n37) );
  DFF_X1 \x_reg[3][7]  ( .D(n215), .CK(clk), .Q(\x[3][7] ), .QN(n1) );
  DFF_X1 \x_reg[0][1]  ( .D(n245), .CK(clk), .Q(\x[0][1] ), .QN(n22) );
  DFF_X1 \x_reg[0][7]  ( .D(n239), .CK(clk), .Q(\x[0][7] ), .QN(n20) );
  DFF_X1 \a_reg[2][3]  ( .D(n355), .CK(clk), .QN(n185) );
  DFF_X1 \a_reg[11][7]  ( .D(n279), .CK(clk), .Q(\a[11][7] ), .QN(n14) );
  INV_X1 U3 ( .A(n104), .ZN(n105) );
  INV_X1 U4 ( .A(n11), .ZN(n13) );
  INV_X2 U5 ( .A(n14), .ZN(n17) );
  INV_X2 U6 ( .A(n185), .ZN(n186) );
  INV_X1 U7 ( .A(n18), .ZN(n19) );
  INV_X2 U8 ( .A(n20), .ZN(n21) );
  INV_X2 U9 ( .A(n22), .ZN(n23) );
  INV_X1 U10 ( .A(n24), .ZN(n25) );
  INV_X1 U11 ( .A(n26), .ZN(n27) );
  INV_X1 U12 ( .A(n28), .ZN(n29) );
  INV_X2 U13 ( .A(n30), .ZN(n31) );
  CLKBUF_X3 U14 ( .A(\x[2][1] ), .Z(n406) );
  INV_X2 U15 ( .A(n1), .ZN(n32) );
  INV_X1 U16 ( .A(n33), .ZN(n34) );
  INV_X1 U17 ( .A(n35), .ZN(n36) );
  INV_X2 U18 ( .A(n37), .ZN(n38) );
  INV_X1 U19 ( .A(n39), .ZN(n41) );
  INV_X2 U20 ( .A(n5), .ZN(n42) );
  INV_X2 U21 ( .A(n43), .ZN(n44) );
  INV_X2 U22 ( .A(n45), .ZN(n46) );
  INV_X2 U23 ( .A(n47), .ZN(n48) );
  INV_X2 U24 ( .A(n49), .ZN(n51) );
  INV_X1 U25 ( .A(n52), .ZN(n53) );
  INV_X1 U26 ( .A(n54), .ZN(n55) );
  CLKBUF_X1 U27 ( .A(n92), .Z(n56) );
  INV_X1 U28 ( .A(n57), .ZN(n58) );
  INV_X2 U29 ( .A(n59), .ZN(n61) );
  INV_X2 U30 ( .A(n62), .ZN(n63) );
  INV_X2 U31 ( .A(n64), .ZN(n65) );
  INV_X1 U32 ( .A(n66), .ZN(n67) );
  INV_X2 U33 ( .A(n68), .ZN(n69) );
  INV_X2 U34 ( .A(n2), .ZN(n72) );
  BUF_X2 U35 ( .A(\x[3][6] ), .Z(n404) );
  INV_X2 U36 ( .A(n3), .ZN(n73) );
  INV_X1 U37 ( .A(n7), .ZN(n74) );
  INV_X2 U38 ( .A(n75), .ZN(n76) );
  INV_X2 U39 ( .A(n77), .ZN(n78) );
  CLKBUF_X1 U40 ( .A(n145), .Z(n79) );
  INV_X2 U41 ( .A(n83), .ZN(n84) );
  INV_X1 U42 ( .A(n85), .ZN(n86) );
  INV_X2 U43 ( .A(n87), .ZN(n88) );
  INV_X2 U44 ( .A(n89), .ZN(n90) );
  INV_X2 U45 ( .A(n91), .ZN(n92) );
  CLKBUF_X1 U46 ( .A(n135), .Z(n93) );
  INV_X2 U47 ( .A(n94), .ZN(n95) );
  INV_X1 U48 ( .A(n97), .ZN(n98) );
  INV_X1 U49 ( .A(n99), .ZN(n100) );
  CLKBUF_X1 U50 ( .A(n105), .Z(n101) );
  INV_X2 U51 ( .A(n102), .ZN(n103) );
  INV_X1 U52 ( .A(n106), .ZN(n107) );
  AND2_X1 U53 ( .A1(N23), .A2(N22), .ZN(n108) );
  AND2_X1 U54 ( .A1(n427), .A2(N23), .ZN(n110) );
  AND2_X1 U55 ( .A1(n193), .A2(n50), .ZN(n111) );
  AND2_X1 U56 ( .A1(n193), .A2(n70), .ZN(n112) );
  AND2_X1 U57 ( .A1(N104), .A2(en_x), .ZN(n113) );
  AND3_X1 U58 ( .A1(n15), .A2(n16), .A3(en_x), .ZN(n114) );
  AND2_X1 U59 ( .A1(n40), .A2(n50), .ZN(n115) );
  AND2_X1 U60 ( .A1(n50), .A2(n119), .ZN(n116) );
  AND2_X1 U61 ( .A1(en_a), .A2(N103), .ZN(n117) );
  AND2_X1 U62 ( .A1(n193), .A2(n60), .ZN(n118) );
  AND3_X1 U63 ( .A1(addr_x[1]), .A2(n16), .A3(en_x), .ZN(n120) );
  AND3_X1 U64 ( .A1(addr_x[0]), .A2(n15), .A3(en_x), .ZN(n121) );
  AND2_X1 U65 ( .A1(n40), .A2(n425), .ZN(n122) );
  AND2_X1 U66 ( .A1(n40), .A2(n60), .ZN(n123) );
  AND2_X1 U67 ( .A1(n40), .A2(n70), .ZN(n124) );
  AND2_X1 U68 ( .A1(n81), .A2(n425), .ZN(n125) );
  AND2_X1 U69 ( .A1(n81), .A2(n50), .ZN(n126) );
  AND2_X1 U70 ( .A1(n81), .A2(n60), .ZN(n127) );
  AND2_X1 U71 ( .A1(n81), .A2(n70), .ZN(n128) );
  AND2_X1 U72 ( .A1(n119), .A2(n425), .ZN(n129) );
  AND2_X1 U73 ( .A1(n60), .A2(n119), .ZN(n130) );
  AND2_X1 U74 ( .A1(n119), .A2(n70), .ZN(n131) );
  AND2_X1 U75 ( .A1(n426), .A2(N22), .ZN(n132) );
  AND2_X1 U76 ( .A1(n426), .A2(n427), .ZN(n133) );
  INV_X2 U77 ( .A(n134), .ZN(n135) );
  INV_X2 U78 ( .A(n136), .ZN(n137) );
  INV_X2 U79 ( .A(n138), .ZN(n139) );
  INV_X2 U80 ( .A(n140), .ZN(n141) );
  INV_X2 U81 ( .A(n142), .ZN(n143) );
  INV_X2 U82 ( .A(n144), .ZN(n145) );
  INV_X2 U83 ( .A(n146), .ZN(n147) );
  INV_X2 U84 ( .A(n148), .ZN(n149) );
  INV_X2 U85 ( .A(n150), .ZN(n151) );
  INV_X2 U86 ( .A(n152), .ZN(n153) );
  INV_X2 U87 ( .A(n154), .ZN(n155) );
  INV_X2 U88 ( .A(n156), .ZN(n157) );
  INV_X2 U89 ( .A(n158), .ZN(n159) );
  INV_X2 U90 ( .A(n160), .ZN(n161) );
  INV_X2 U91 ( .A(n162), .ZN(n163) );
  INV_X2 U92 ( .A(n164), .ZN(n165) );
  INV_X2 U93 ( .A(n166), .ZN(n167) );
  CLKBUF_X1 U94 ( .A(n41), .Z(n168) );
  INV_X2 U95 ( .A(n169), .ZN(n170) );
  INV_X2 U96 ( .A(n171), .ZN(n172) );
  INV_X2 U97 ( .A(n173), .ZN(n174) );
  INV_X1 U98 ( .A(n175), .ZN(n176) );
  INV_X2 U99 ( .A(n177), .ZN(n178) );
  INV_X1 U100 ( .A(n179), .ZN(n180) );
  INV_X1 U101 ( .A(n181), .ZN(n182) );
  INV_X2 U102 ( .A(n183), .ZN(n184) );
  INV_X2 U103 ( .A(n187), .ZN(n188) );
  INV_X2 U104 ( .A(n189), .ZN(n190) );
  INV_X2 U105 ( .A(n191), .ZN(n192) );
  INV_X1 U106 ( .A(n194), .ZN(n195) );
  INV_X2 U107 ( .A(n196), .ZN(n197) );
  INV_X2 U108 ( .A(n198), .ZN(n199) );
  INV_X2 U109 ( .A(n200), .ZN(n201) );
  INV_X2 U110 ( .A(n202), .ZN(n203) );
  INV_X1 U111 ( .A(n213), .ZN(n428) );
  OAI21_X1 U112 ( .B1(n50), .B2(n60), .A(n429), .ZN(n213) );
  NOR2_X1 U113 ( .A1(n15), .A2(n16), .ZN(N104) );
  NOR3_X1 U114 ( .A1(n10), .A2(n9), .A3(n211), .ZN(N103) );
  NOR2_X1 U115 ( .A1(n12), .A2(addr_a[0]), .ZN(n50) );
  AOI21_X1 U116 ( .B1(n429), .B2(n12), .A(N87), .ZN(n208) );
  NOR2_X1 U117 ( .A1(addr_a[0]), .A2(addr_a[1]), .ZN(n70) );
  OAI22_X1 U118 ( .A1(n208), .A2(n9), .B1(clr_addr_a), .B2(n209), .ZN(N90) );
  AOI22_X1 U119 ( .A1(n210), .A2(n425), .B1(addr_a[3]), .B2(n10), .ZN(n209) );
  NOR2_X1 U120 ( .A1(addr_a[3]), .A2(n10), .ZN(n210) );
  OAI22_X1 U121 ( .A1(n208), .A2(n10), .B1(n211), .B2(n212), .ZN(N89) );
  NAND2_X1 U122 ( .A1(n10), .A2(n429), .ZN(n212) );
  NOR2_X1 U123 ( .A1(addr_a[0]), .A2(clr_addr_a), .ZN(N87) );
  AND2_X1 U124 ( .A1(addr_a[0]), .A2(n12), .ZN(n60) );
  NAND2_X1 U125 ( .A1(addr_a[1]), .A2(addr_a[0]), .ZN(n211) );
  INV_X1 U126 ( .A(clr_addr_a), .ZN(n429) );
  AND2_X1 U127 ( .A1(n109), .A2(n10), .ZN(n119) );
  AND2_X1 U128 ( .A1(n71), .A2(n10), .ZN(n40) );
  AND2_X1 U129 ( .A1(n109), .A2(addr_a[2]), .ZN(n81) );
  BUF_X1 U130 ( .A(\x[1][0] ), .Z(n408) );
  NOR2_X1 U131 ( .A1(clr_addr_y), .A2(n214), .ZN(N100) );
  XNOR2_X1 U132 ( .A(N23), .B(N22), .ZN(n214) );
  NOR2_X1 U133 ( .A1(clr_addr_y), .A2(N22), .ZN(N99) );
  NOR2_X1 U134 ( .A1(clr_addr_x), .A2(n207), .ZN(N95) );
  NOR2_X1 U135 ( .A1(clr_addr_x), .A2(addr_x[0]), .ZN(N94) );
  AND2_X1 U136 ( .A1(addr_a[2]), .A2(n71), .ZN(n193) );
  AND2_X1 U137 ( .A1(N22), .A2(N23), .ZN(N105) );
  AND2_X1 U138 ( .A1(en_a), .A2(addr_a[3]), .ZN(n71) );
  AND2_X1 U139 ( .A1(en_a), .A2(n9), .ZN(n109) );
  MUX2_X1 U140 ( .A(\y[2][0] ), .B(\y[3][0] ), .S(N22), .Z(n204) );
  MUX2_X1 U141 ( .A(\y[0][0] ), .B(\y[1][0] ), .S(N22), .Z(n205) );
  MUX2_X1 U142 ( .A(n205), .B(n204), .S(N23), .Z(N81) );
  MUX2_X1 U143 ( .A(\y[2][1] ), .B(\y[3][1] ), .S(N22), .Z(n206) );
  MUX2_X1 U144 ( .A(\y[0][1] ), .B(\y[1][1] ), .S(N22), .Z(n375) );
  MUX2_X1 U145 ( .A(n375), .B(n206), .S(N23), .Z(N80) );
  MUX2_X1 U146 ( .A(\y[2][2] ), .B(\y[3][2] ), .S(N22), .Z(n376) );
  MUX2_X1 U147 ( .A(\y[0][2] ), .B(\y[1][2] ), .S(N22), .Z(n377) );
  MUX2_X1 U148 ( .A(n377), .B(n376), .S(N23), .Z(N79) );
  MUX2_X1 U149 ( .A(\y[2][3] ), .B(\y[3][3] ), .S(N22), .Z(n378) );
  MUX2_X1 U150 ( .A(\y[0][3] ), .B(\y[1][3] ), .S(N22), .Z(n379) );
  MUX2_X1 U151 ( .A(\y[2][4] ), .B(\y[3][4] ), .S(N22), .Z(n380) );
  MUX2_X1 U152 ( .A(\y[0][4] ), .B(\y[1][4] ), .S(N22), .Z(n381) );
  MUX2_X1 U153 ( .A(n381), .B(n380), .S(N23), .Z(N77) );
  MUX2_X1 U154 ( .A(\y[2][5] ), .B(\y[3][5] ), .S(N22), .Z(n382) );
  MUX2_X1 U155 ( .A(\y[0][5] ), .B(\y[1][5] ), .S(N22), .Z(n383) );
  MUX2_X1 U156 ( .A(n383), .B(n382), .S(N23), .Z(N76) );
  MUX2_X1 U157 ( .A(\y[2][6] ), .B(\y[3][6] ), .S(N22), .Z(n384) );
  MUX2_X1 U158 ( .A(\y[0][6] ), .B(\y[1][6] ), .S(N22), .Z(n385) );
  MUX2_X1 U159 ( .A(n385), .B(n384), .S(N23), .Z(N75) );
  MUX2_X1 U160 ( .A(\y[2][7] ), .B(\y[3][7] ), .S(N22), .Z(n386) );
  MUX2_X1 U161 ( .A(\y[0][7] ), .B(\y[1][7] ), .S(N22), .Z(n387) );
  MUX2_X1 U162 ( .A(n387), .B(n386), .S(N23), .Z(N74) );
  MUX2_X1 U163 ( .A(\y[2][8] ), .B(\y[3][8] ), .S(N22), .Z(n388) );
  MUX2_X1 U164 ( .A(\y[0][8] ), .B(\y[1][8] ), .S(N22), .Z(n389) );
  MUX2_X1 U165 ( .A(n389), .B(n388), .S(N23), .Z(N73) );
  NAND2_X1 U166 ( .A1(n390), .A2(n391), .ZN(N72) );
  AOI22_X1 U167 ( .A1(\y[2][9] ), .A2(n110), .B1(\y[0][9] ), .B2(n133), .ZN(
        n391) );
  AOI22_X1 U168 ( .A1(\y[3][9] ), .A2(n108), .B1(\y[1][9] ), .B2(n132), .ZN(
        n390) );
  NAND2_X1 U169 ( .A1(n392), .A2(n393), .ZN(N71) );
  AOI22_X1 U170 ( .A1(\y[2][10] ), .A2(n110), .B1(\y[0][10] ), .B2(n133), .ZN(
        n393) );
  AOI22_X1 U171 ( .A1(\y[3][10] ), .A2(n108), .B1(\y[1][10] ), .B2(n132), .ZN(
        n392) );
  NAND2_X1 U172 ( .A1(n394), .A2(n395), .ZN(N70) );
  AOI22_X1 U173 ( .A1(\y[2][11] ), .A2(n110), .B1(\y[0][11] ), .B2(n133), .ZN(
        n395) );
  AOI22_X1 U174 ( .A1(\y[3][11] ), .A2(n108), .B1(\y[1][11] ), .B2(n132), .ZN(
        n394) );
  NAND2_X1 U175 ( .A1(n396), .A2(n397), .ZN(N69) );
  AOI22_X1 U176 ( .A1(\y[2][12] ), .A2(n110), .B1(\y[0][12] ), .B2(n133), .ZN(
        n397) );
  AOI22_X1 U177 ( .A1(\y[3][12] ), .A2(n108), .B1(\y[1][12] ), .B2(n132), .ZN(
        n396) );
  NAND2_X1 U178 ( .A1(n398), .A2(n399), .ZN(N68) );
  AOI22_X1 U179 ( .A1(\y[2][13] ), .A2(n110), .B1(\y[0][13] ), .B2(n133), .ZN(
        n399) );
  AOI22_X1 U180 ( .A1(\y[3][13] ), .A2(n108), .B1(\y[1][13] ), .B2(n132), .ZN(
        n398) );
  NAND2_X1 U181 ( .A1(n400), .A2(n401), .ZN(N67) );
  AOI22_X1 U182 ( .A1(\y[2][14] ), .A2(n110), .B1(\y[0][14] ), .B2(n133), .ZN(
        n401) );
  AOI22_X1 U183 ( .A1(\y[3][14] ), .A2(n108), .B1(\y[1][14] ), .B2(n132), .ZN(
        n400) );
  NAND2_X1 U184 ( .A1(n402), .A2(n403), .ZN(N66) );
  AOI22_X1 U185 ( .A1(\y[2][15] ), .A2(n110), .B1(\y[0][15] ), .B2(n133), .ZN(
        n403) );
  AOI22_X1 U186 ( .A1(\y[3][15] ), .A2(n108), .B1(\y[1][15] ), .B2(n132), .ZN(
        n402) );
  BUF_X4 U187 ( .A(\x[2][2] ), .Z(n405) );
  BUF_X4 U188 ( .A(\x[3][5] ), .Z(n407) );
  MUX2_X1 U189 ( .A(\a[15][7] ), .B(data_in[7]), .S(n117), .Z(n247) );
  MUX2_X1 U190 ( .A(\a[15][6] ), .B(data_in[6]), .S(n117), .Z(n248) );
  MUX2_X1 U191 ( .A(\a[15][5] ), .B(data_in[5]), .S(n117), .Z(n249) );
  MUX2_X1 U192 ( .A(\a[15][4] ), .B(data_in[4]), .S(n117), .Z(n250) );
  MUX2_X1 U193 ( .A(n80), .B(data_in[3]), .S(n117), .Z(n251) );
  MUX2_X1 U194 ( .A(\a[15][2] ), .B(data_in[2]), .S(n117), .Z(n252) );
  MUX2_X1 U195 ( .A(\a[15][1] ), .B(data_in[1]), .S(n117), .Z(n253) );
  MUX2_X1 U196 ( .A(\a[15][0] ), .B(data_in[0]), .S(n117), .Z(n254) );
  MUX2_X1 U197 ( .A(n36), .B(data_in[7]), .S(n111), .Z(n255) );
  MUX2_X1 U198 ( .A(\a[14][6] ), .B(data_in[6]), .S(n111), .Z(n256) );
  MUX2_X1 U199 ( .A(n55), .B(data_in[5]), .S(n111), .Z(n257) );
  MUX2_X1 U200 ( .A(\a[14][4] ), .B(data_in[4]), .S(n111), .Z(n258) );
  MUX2_X1 U201 ( .A(\a[14][3] ), .B(data_in[3]), .S(n111), .Z(n259) );
  MUX2_X1 U202 ( .A(\a[14][2] ), .B(data_in[2]), .S(n111), .Z(n260) );
  MUX2_X1 U203 ( .A(n29), .B(data_in[1]), .S(n111), .Z(n261) );
  MUX2_X1 U204 ( .A(\a[14][0] ), .B(data_in[0]), .S(n111), .Z(n262) );
  MUX2_X1 U205 ( .A(n82), .B(data_in[7]), .S(n118), .Z(n263) );
  MUX2_X1 U206 ( .A(\a[13][6] ), .B(data_in[6]), .S(n118), .Z(n264) );
  MUX2_X1 U207 ( .A(\a[13][5] ), .B(data_in[5]), .S(n118), .Z(n265) );
  MUX2_X1 U208 ( .A(\a[13][4] ), .B(data_in[4]), .S(n118), .Z(n266) );
  MUX2_X1 U209 ( .A(\a[13][3] ), .B(data_in[3]), .S(n118), .Z(n267) );
  MUX2_X1 U210 ( .A(\a[13][2] ), .B(data_in[2]), .S(n118), .Z(n268) );
  MUX2_X1 U211 ( .A(n25), .B(data_in[1]), .S(n118), .Z(n269) );
  MUX2_X1 U212 ( .A(\a[13][0] ), .B(data_in[0]), .S(n118), .Z(n270) );
  MUX2_X1 U213 ( .A(n95), .B(data_in[7]), .S(n112), .Z(n271) );
  MUX2_X1 U214 ( .A(\a[12][6] ), .B(data_in[6]), .S(n112), .Z(n272) );
  MUX2_X1 U215 ( .A(\a[12][5] ), .B(data_in[5]), .S(n112), .Z(n273) );
  MUX2_X1 U216 ( .A(\a[12][4] ), .B(data_in[4]), .S(n112), .Z(n274) );
  MUX2_X1 U217 ( .A(\a[12][3] ), .B(data_in[3]), .S(n112), .Z(n275) );
  MUX2_X1 U218 ( .A(\a[12][2] ), .B(data_in[2]), .S(n112), .Z(n276) );
  MUX2_X1 U219 ( .A(\a[12][1] ), .B(data_in[1]), .S(n112), .Z(n277) );
  MUX2_X1 U220 ( .A(\a[12][0] ), .B(data_in[0]), .S(n112), .Z(n278) );
  INV_X1 U221 ( .A(data_in[7]), .ZN(n409) );
  MUX2_X1 U222 ( .A(n1), .B(n409), .S(n113), .Z(n410) );
  INV_X1 U223 ( .A(n410), .ZN(n215) );
  INV_X1 U224 ( .A(data_in[6]), .ZN(n411) );
  MUX2_X1 U225 ( .A(n2), .B(n411), .S(n113), .Z(n412) );
  INV_X1 U226 ( .A(n412), .ZN(n216) );
  INV_X1 U227 ( .A(data_in[5]), .ZN(n413) );
  MUX2_X1 U228 ( .A(n3), .B(n413), .S(n113), .Z(n414) );
  INV_X1 U229 ( .A(n414), .ZN(n217) );
  INV_X1 U230 ( .A(data_in[4]), .ZN(n415) );
  MUX2_X1 U231 ( .A(n4), .B(n415), .S(n113), .Z(n416) );
  INV_X1 U232 ( .A(n416), .ZN(n218) );
  INV_X1 U233 ( .A(data_in[3]), .ZN(n417) );
  MUX2_X1 U234 ( .A(n5), .B(n417), .S(n113), .Z(n418) );
  INV_X1 U235 ( .A(n418), .ZN(n219) );
  INV_X1 U236 ( .A(data_in[2]), .ZN(n419) );
  MUX2_X1 U237 ( .A(n6), .B(n419), .S(n113), .Z(n420) );
  INV_X1 U238 ( .A(n420), .ZN(n220) );
  INV_X1 U239 ( .A(data_in[1]), .ZN(n421) );
  MUX2_X1 U240 ( .A(n7), .B(n421), .S(n113), .Z(n422) );
  INV_X1 U241 ( .A(n422), .ZN(n221) );
  INV_X1 U242 ( .A(data_in[0]), .ZN(n423) );
  MUX2_X1 U243 ( .A(n8), .B(n423), .S(n113), .Z(n424) );
  INV_X1 U244 ( .A(n424), .ZN(n222) );
  MUX2_X1 U245 ( .A(\x[2][7] ), .B(data_in[7]), .S(n120), .Z(n223) );
  MUX2_X1 U246 ( .A(n38), .B(data_in[6]), .S(n120), .Z(n224) );
  MUX2_X1 U247 ( .A(n44), .B(data_in[5]), .S(n120), .Z(n225) );
  MUX2_X1 U248 ( .A(n65), .B(data_in[4]), .S(n120), .Z(n226) );
  MUX2_X1 U249 ( .A(n61), .B(data_in[3]), .S(n120), .Z(n227) );
  MUX2_X1 U250 ( .A(n405), .B(data_in[2]), .S(n120), .Z(n228) );
  MUX2_X1 U251 ( .A(n31), .B(data_in[1]), .S(n120), .Z(n229) );
  MUX2_X1 U252 ( .A(n100), .B(data_in[0]), .S(n120), .Z(n230) );
  MUX2_X1 U253 ( .A(\x[1][7] ), .B(data_in[7]), .S(n121), .Z(n231) );
  MUX2_X1 U254 ( .A(n46), .B(data_in[6]), .S(n121), .Z(n232) );
  MUX2_X1 U255 ( .A(n48), .B(data_in[5]), .S(n121), .Z(n233) );
  MUX2_X1 U256 ( .A(\x[1][4] ), .B(data_in[4]), .S(n121), .Z(n234) );
  MUX2_X1 U257 ( .A(\x[1][3] ), .B(data_in[3]), .S(n121), .Z(n235) );
  MUX2_X1 U258 ( .A(\x[1][2] ), .B(data_in[2]), .S(n121), .Z(n236) );
  MUX2_X1 U259 ( .A(n188), .B(data_in[1]), .S(n121), .Z(n237) );
  MUX2_X1 U260 ( .A(n408), .B(data_in[0]), .S(n121), .Z(n238) );
  MUX2_X1 U261 ( .A(n21), .B(data_in[7]), .S(n114), .Z(n239) );
  MUX2_X1 U262 ( .A(n170), .B(data_in[6]), .S(n114), .Z(n240) );
  MUX2_X1 U263 ( .A(n178), .B(data_in[5]), .S(n114), .Z(n241) );
  MUX2_X1 U264 ( .A(\x[0][4] ), .B(data_in[4]), .S(n114), .Z(n242) );
  MUX2_X1 U265 ( .A(\x[0][3] ), .B(data_in[3]), .S(n114), .Z(n243) );
  MUX2_X1 U266 ( .A(\x[0][2] ), .B(data_in[2]), .S(n114), .Z(n244) );
  MUX2_X1 U267 ( .A(n23), .B(data_in[1]), .S(n114), .Z(n245) );
  MUX2_X1 U268 ( .A(\x[0][0] ), .B(data_in[0]), .S(n114), .Z(n246) );
  INV_X1 U269 ( .A(n211), .ZN(n425) );
  MUX2_X1 U270 ( .A(\a[11][7] ), .B(data_in[7]), .S(n122), .Z(n279) );
  MUX2_X1 U271 ( .A(\a[11][6] ), .B(data_in[6]), .S(n122), .Z(n280) );
  MUX2_X1 U272 ( .A(n86), .B(data_in[5]), .S(n122), .Z(n281) );
  MUX2_X1 U273 ( .A(\a[11][4] ), .B(data_in[4]), .S(n122), .Z(n282) );
  MUX2_X1 U274 ( .A(\a[11][3] ), .B(data_in[3]), .S(n122), .Z(n283) );
  MUX2_X1 U275 ( .A(\a[11][2] ), .B(data_in[2]), .S(n122), .Z(n284) );
  MUX2_X1 U276 ( .A(\a[11][1] ), .B(data_in[1]), .S(n122), .Z(n285) );
  MUX2_X1 U277 ( .A(\a[11][0] ), .B(data_in[0]), .S(n122), .Z(n286) );
  MUX2_X1 U278 ( .A(n79), .B(data_in[7]), .S(n115), .Z(n287) );
  MUX2_X1 U279 ( .A(\a[10][6] ), .B(data_in[6]), .S(n115), .Z(n288) );
  MUX2_X1 U280 ( .A(n98), .B(data_in[5]), .S(n115), .Z(n289) );
  MUX2_X1 U281 ( .A(\a[10][4] ), .B(data_in[4]), .S(n115), .Z(n290) );
  MUX2_X1 U282 ( .A(n93), .B(data_in[3]), .S(n115), .Z(n291) );
  MUX2_X1 U283 ( .A(\a[10][2] ), .B(data_in[2]), .S(n115), .Z(n292) );
  MUX2_X1 U284 ( .A(n19), .B(data_in[1]), .S(n115), .Z(n293) );
  MUX2_X1 U285 ( .A(\a[10][0] ), .B(data_in[0]), .S(n115), .Z(n294) );
  MUX2_X1 U286 ( .A(n96), .B(data_in[7]), .S(n123), .Z(n295) );
  MUX2_X1 U287 ( .A(\a[9][6] ), .B(data_in[6]), .S(n123), .Z(n296) );
  MUX2_X1 U288 ( .A(\a[9][5] ), .B(data_in[5]), .S(n123), .Z(n297) );
  MUX2_X1 U289 ( .A(\a[9][4] ), .B(data_in[4]), .S(n123), .Z(n298) );
  MUX2_X1 U290 ( .A(\a[9][3] ), .B(data_in[3]), .S(n123), .Z(n299) );
  MUX2_X1 U291 ( .A(\a[9][2] ), .B(data_in[2]), .S(n123), .Z(n300) );
  MUX2_X1 U292 ( .A(n13), .B(data_in[1]), .S(n123), .Z(n301) );
  MUX2_X1 U293 ( .A(\a[9][0] ), .B(data_in[0]), .S(n123), .Z(n302) );
  MUX2_X1 U294 ( .A(\a[8][7] ), .B(data_in[7]), .S(n124), .Z(n303) );
  MUX2_X1 U295 ( .A(\a[8][6] ), .B(data_in[6]), .S(n124), .Z(n304) );
  MUX2_X1 U296 ( .A(\a[8][5] ), .B(data_in[5]), .S(n124), .Z(n305) );
  MUX2_X1 U297 ( .A(\a[8][4] ), .B(data_in[4]), .S(n124), .Z(n306) );
  MUX2_X1 U298 ( .A(\a[8][3] ), .B(data_in[3]), .S(n124), .Z(n307) );
  MUX2_X1 U299 ( .A(\a[8][2] ), .B(data_in[2]), .S(n124), .Z(n308) );
  MUX2_X1 U300 ( .A(\a[8][1] ), .B(data_in[1]), .S(n124), .Z(n309) );
  MUX2_X1 U301 ( .A(\a[8][0] ), .B(data_in[0]), .S(n124), .Z(n310) );
  MUX2_X1 U302 ( .A(n165), .B(data_in[7]), .S(n125), .Z(n311) );
  MUX2_X1 U303 ( .A(\a[7][6] ), .B(data_in[6]), .S(n125), .Z(n312) );
  MUX2_X1 U304 ( .A(n195), .B(data_in[5]), .S(n125), .Z(n313) );
  MUX2_X1 U305 ( .A(\a[7][4] ), .B(data_in[4]), .S(n125), .Z(n314) );
  MUX2_X1 U306 ( .A(\a[7][3] ), .B(data_in[3]), .S(n125), .Z(n315) );
  MUX2_X1 U307 ( .A(\a[7][2] ), .B(data_in[2]), .S(n125), .Z(n316) );
  MUX2_X1 U308 ( .A(n101), .B(data_in[1]), .S(n125), .Z(n317) );
  MUX2_X1 U309 ( .A(\a[7][0] ), .B(data_in[0]), .S(n125), .Z(n318) );
  MUX2_X1 U310 ( .A(\a[6][7] ), .B(data_in[7]), .S(n126), .Z(n319) );
  MUX2_X1 U311 ( .A(\a[6][6] ), .B(data_in[6]), .S(n126), .Z(n320) );
  MUX2_X1 U312 ( .A(n27), .B(data_in[5]), .S(n126), .Z(n321) );
  MUX2_X1 U313 ( .A(\a[6][4] ), .B(data_in[4]), .S(n126), .Z(n322) );
  MUX2_X1 U314 ( .A(n180), .B(data_in[3]), .S(n126), .Z(n323) );
  MUX2_X1 U315 ( .A(\a[6][2] ), .B(data_in[2]), .S(n126), .Z(n324) );
  MUX2_X1 U316 ( .A(\a[6][1] ), .B(data_in[1]), .S(n126), .Z(n325) );
  MUX2_X1 U317 ( .A(\a[6][0] ), .B(data_in[0]), .S(n126), .Z(n326) );
  MUX2_X1 U318 ( .A(n67), .B(data_in[7]), .S(n127), .Z(n327) );
  MUX2_X1 U319 ( .A(\a[5][6] ), .B(data_in[6]), .S(n127), .Z(n328) );
  MUX2_X1 U320 ( .A(\a[5][5] ), .B(data_in[5]), .S(n127), .Z(n329) );
  MUX2_X1 U321 ( .A(\a[5][4] ), .B(data_in[4]), .S(n127), .Z(n330) );
  MUX2_X1 U322 ( .A(n56), .B(data_in[3]), .S(n127), .Z(n331) );
  MUX2_X1 U323 ( .A(\a[5][2] ), .B(data_in[2]), .S(n127), .Z(n332) );
  MUX2_X1 U324 ( .A(\a[5][1] ), .B(data_in[1]), .S(n127), .Z(n333) );
  MUX2_X1 U325 ( .A(\a[5][0] ), .B(data_in[0]), .S(n127), .Z(n334) );
  MUX2_X1 U326 ( .A(\a[4][7] ), .B(data_in[7]), .S(n128), .Z(n335) );
  MUX2_X1 U327 ( .A(\a[4][6] ), .B(data_in[6]), .S(n128), .Z(n336) );
  MUX2_X1 U328 ( .A(\a[4][5] ), .B(data_in[5]), .S(n128), .Z(n337) );
  MUX2_X1 U329 ( .A(\a[4][4] ), .B(data_in[4]), .S(n128), .Z(n338) );
  MUX2_X1 U330 ( .A(n203), .B(data_in[3]), .S(n128), .Z(n339) );
  MUX2_X1 U331 ( .A(\a[4][2] ), .B(data_in[2]), .S(n128), .Z(n340) );
  MUX2_X1 U332 ( .A(\a[4][1] ), .B(data_in[1]), .S(n128), .Z(n341) );
  MUX2_X1 U333 ( .A(\a[4][0] ), .B(data_in[0]), .S(n128), .Z(n342) );
  MUX2_X1 U334 ( .A(\a[3][7] ), .B(data_in[7]), .S(n129), .Z(n343) );
  MUX2_X1 U335 ( .A(\a[3][6] ), .B(data_in[6]), .S(n129), .Z(n344) );
  MUX2_X1 U336 ( .A(n168), .B(data_in[5]), .S(n129), .Z(n345) );
  MUX2_X1 U337 ( .A(\a[3][4] ), .B(data_in[4]), .S(n129), .Z(n346) );
  MUX2_X1 U338 ( .A(n182), .B(data_in[3]), .S(n129), .Z(n347) );
  MUX2_X1 U339 ( .A(\a[3][2] ), .B(data_in[2]), .S(n129), .Z(n348) );
  MUX2_X1 U340 ( .A(n58), .B(data_in[1]), .S(n129), .Z(n349) );
  MUX2_X1 U341 ( .A(\a[3][0] ), .B(data_in[0]), .S(n129), .Z(n350) );
  MUX2_X1 U342 ( .A(\a[2][7] ), .B(data_in[7]), .S(n116), .Z(n351) );
  MUX2_X1 U343 ( .A(\a[2][6] ), .B(data_in[6]), .S(n116), .Z(n352) );
  MUX2_X1 U344 ( .A(\a[2][5] ), .B(data_in[5]), .S(n116), .Z(n353) );
  MUX2_X1 U345 ( .A(\a[2][4] ), .B(data_in[4]), .S(n116), .Z(n354) );
  MUX2_X1 U346 ( .A(n186), .B(data_in[3]), .S(n116), .Z(n355) );
  MUX2_X1 U347 ( .A(n53), .B(data_in[2]), .S(n116), .Z(n356) );
  MUX2_X1 U348 ( .A(n34), .B(data_in[1]), .S(n116), .Z(n357) );
  MUX2_X1 U349 ( .A(\a[2][0] ), .B(data_in[0]), .S(n116), .Z(n358) );
  MUX2_X1 U350 ( .A(\a[1][7] ), .B(data_in[7]), .S(n130), .Z(n359) );
  MUX2_X1 U351 ( .A(\a[1][6] ), .B(data_in[6]), .S(n130), .Z(n360) );
  MUX2_X1 U352 ( .A(\a[1][5] ), .B(data_in[5]), .S(n130), .Z(n361) );
  MUX2_X1 U353 ( .A(\a[1][4] ), .B(data_in[4]), .S(n130), .Z(n362) );
  MUX2_X1 U354 ( .A(\a[1][3] ), .B(data_in[3]), .S(n130), .Z(n363) );
  MUX2_X1 U355 ( .A(\a[1][2] ), .B(data_in[2]), .S(n130), .Z(n364) );
  MUX2_X1 U356 ( .A(\a[1][1] ), .B(data_in[1]), .S(n130), .Z(n365) );
  MUX2_X1 U357 ( .A(\a[1][0] ), .B(data_in[0]), .S(n130), .Z(n366) );
  MUX2_X1 U358 ( .A(\a[0][7] ), .B(data_in[7]), .S(n131), .Z(n367) );
  MUX2_X1 U359 ( .A(\a[0][6] ), .B(data_in[6]), .S(n131), .Z(n368) );
  MUX2_X1 U360 ( .A(\a[0][5] ), .B(data_in[5]), .S(n131), .Z(n369) );
  MUX2_X1 U361 ( .A(n107), .B(data_in[4]), .S(n131), .Z(n370) );
  MUX2_X1 U362 ( .A(n176), .B(data_in[3]), .S(n131), .Z(n371) );
  MUX2_X1 U363 ( .A(\a[0][2] ), .B(data_in[2]), .S(n131), .Z(n372) );
  MUX2_X1 U364 ( .A(\a[0][1] ), .B(data_in[1]), .S(n131), .Z(n373) );
  MUX2_X1 U365 ( .A(\a[0][0] ), .B(data_in[0]), .S(n131), .Z(n374) );
endmodule


module control ( clk, reset, start, done, en_a, en_x, en_y, clr_addr_a, 
        clr_addr_x, clr_addr_y, of_a, of_x, of_y );
  input clk, reset, start, of_a, of_x, of_y;
  output done, en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y;
  wire   \out_state[0] , n7, n9, n11, n12, n13, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n1,
         n2, n3, n4, n5, n6, n8, n10, n14, n15, n16;
  wire   [1:0] in_state;

  DFF_X1 done_reg ( .D(n6), .CK(clk), .Q(done) );
  DFF_X1 en_a_reg ( .D(n47), .CK(clk), .Q(en_a) );
  DFF_X1 en_x_reg ( .D(n46), .CK(clk), .Q(en_x) );
  DFF_X1 en_y_reg ( .D(n8), .CK(clk), .Q(en_y) );
  DFF_X1 clr_addr_y_reg ( .D(n43), .CK(clk), .Q(clr_addr_y) );
  NAND3_X1 U46 ( .A1(n3), .A2(n15), .A3(n23), .ZN(n28) );
  NAND3_X1 U47 ( .A1(n38), .A2(n15), .A3(n23), .ZN(n39) );
  NAND3_X1 U48 ( .A1(n38), .A2(n15), .A3(n41), .ZN(n40) );
  DFF_X1 \out_state_reg[0]  ( .D(n48), .CK(clk), .Q(\out_state[0] ), .QN(n11)
         );
  DFF_X1 clr_addr_a_reg ( .D(n45), .CK(clk), .Q(clr_addr_a), .QN(n12) );
  DFF_X1 clr_addr_x_reg ( .D(n44), .CK(clk), .Q(clr_addr_x), .QN(n13) );
  DFF_X1 \in_state_reg[1]  ( .D(n49), .CK(clk), .Q(in_state[1]), .QN(n7) );
  DFF_X1 \in_state_reg[0]  ( .D(n50), .CK(clk), .Q(in_state[0]), .QN(n9) );
  INV_X1 U3 ( .A(n19), .ZN(n3) );
  INV_X1 U4 ( .A(n21), .ZN(n1) );
  OAI21_X1 U5 ( .B1(n16), .B2(n33), .A(n19), .ZN(n38) );
  OAI21_X1 U6 ( .B1(n31), .B2(n16), .A(n32), .ZN(n21) );
  AOI21_X1 U7 ( .B1(n4), .B2(of_x), .A(n2), .ZN(n31) );
  INV_X1 U8 ( .A(n42), .ZN(n4) );
  INV_X1 U9 ( .A(n33), .ZN(n2) );
  AOI21_X1 U10 ( .B1(of_x), .B2(n4), .A(n5), .ZN(n19) );
  INV_X1 U11 ( .A(n32), .ZN(n5) );
  NOR2_X1 U12 ( .A1(n9), .A2(in_state[1]), .ZN(n23) );
  NOR2_X1 U13 ( .A1(n18), .A2(in_state[0]), .ZN(n25) );
  AOI21_X1 U14 ( .B1(n23), .B2(of_a), .A(reset), .ZN(n32) );
  OAI22_X1 U15 ( .A1(n3), .A2(n13), .B1(n19), .B2(n20), .ZN(n44) );
  NOR2_X1 U16 ( .A1(n4), .A2(reset), .ZN(n20) );
  OAI22_X1 U17 ( .A1(n21), .A2(n12), .B1(n1), .B2(n22), .ZN(n45) );
  NOR2_X1 U18 ( .A1(n23), .A2(reset), .ZN(n22) );
  NAND2_X1 U19 ( .A1(n9), .A2(n7), .ZN(n33) );
  AOI21_X1 U20 ( .B1(n36), .B2(n37), .A(reset), .ZN(n48) );
  NAND2_X1 U21 ( .A1(n14), .A2(\out_state[0] ), .ZN(n37) );
  NAND2_X1 U22 ( .A1(n25), .A2(n11), .ZN(n36) );
  OAI21_X1 U23 ( .B1(n9), .B2(n38), .A(n40), .ZN(n50) );
  OAI21_X1 U24 ( .B1(n42), .B2(n16), .A(n33), .ZN(n41) );
  NAND2_X1 U25 ( .A1(of_x), .A2(in_state[1]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(in_state[1]), .A2(n9), .ZN(n42) );
  OAI21_X1 U27 ( .B1(n7), .B2(n38), .A(n39), .ZN(n49) );
  INV_X1 U28 ( .A(n26), .ZN(n10) );
  OAI21_X1 U29 ( .B1(n11), .B2(n14), .A(n15), .ZN(n26) );
  INV_X1 U30 ( .A(of_y), .ZN(n14) );
  NAND2_X1 U31 ( .A1(n29), .A2(n30), .ZN(n47) );
  OAI211_X1 U32 ( .C1(n2), .C2(n4), .A(n21), .B(n15), .ZN(n30) );
  NAND2_X1 U33 ( .A1(en_a), .A2(n1), .ZN(n29) );
  NAND2_X1 U34 ( .A1(n27), .A2(n28), .ZN(n46) );
  NAND2_X1 U35 ( .A1(en_x), .A2(n19), .ZN(n27) );
  NAND2_X1 U36 ( .A1(n10), .A2(n17), .ZN(n43) );
  OAI21_X1 U37 ( .B1(in_state[0]), .B2(n18), .A(clr_addr_y), .ZN(n17) );
  INV_X1 U38 ( .A(n34), .ZN(n6) );
  OAI211_X1 U39 ( .C1(done), .C2(n25), .A(n11), .B(n15), .ZN(n34) );
  INV_X1 U40 ( .A(n24), .ZN(n8) );
  OAI21_X1 U41 ( .B1(n25), .B2(en_y), .A(n10), .ZN(n24) );
  INV_X1 U42 ( .A(reset), .ZN(n15) );
  INV_X1 U43 ( .A(start), .ZN(n16) );
endmodule


module mvm4_part3 ( clk, reset, start, done, data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, start;
  output done;
  wire   en_a, en_x, en_y, clr_addr_a, clr_addr_x, clr_addr_y, of_a, of_x,
         of_y;

  data_path_MAT_SCALE4_INPUT_WIDTH8_OUTPUT_WIDTH16 datapath ( .clk(clk), 
        .en_a(en_a), .en_x(en_x), .en_y(en_y), .clr_addr_a(clr_addr_a), 
        .clr_addr_x(clr_addr_x), .clr_addr_y(clr_addr_y), .of_a(of_a), .of_x(
        of_x), .of_y(of_y), .data_in(data_in), .data_out(data_out) );
  control ctrl ( .clk(clk), .reset(reset), .start(start), .done(done), .en_a(
        en_a), .en_x(en_x), .en_y(en_y), .clr_addr_a(clr_addr_a), .clr_addr_x(
        clr_addr_x), .clr_addr_y(clr_addr_y), .of_a(of_a), .of_x(of_x), .of_y(
        of_y) );
endmodule

